 /*                                                                      
 Copyright 2018-2020 Nuclei System Technology, Inc.                
                                                                         
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
  Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.                                          
 */                                                                      
                                                                         
                                                                         
                                                                         

module sirv_aon(
  input   clock,
  input   reset,
  input   erst,
  input   test_mode,
  output  io_interrupts_0_0,
  output  io_interrupts_0_1,
  output  io_in_0_a_ready,
  input   io_in_0_a_valid,
  input  [2:0] io_in_0_a_bits_opcode,
  input  [2:0] io_in_0_a_bits_param,
  input  [2:0] io_in_0_a_bits_size,
  input  [4:0] io_in_0_a_bits_source,
  input  [28:0] io_in_0_a_bits_address,
  input  [3:0] io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input   io_in_0_b_ready,
  output  io_in_0_b_valid,
  output [2:0] io_in_0_b_bits_opcode,
  output [1:0] io_in_0_b_bits_param,
  output [2:0] io_in_0_b_bits_size,
  output [4:0] io_in_0_b_bits_source,
  output [28:0] io_in_0_b_bits_address,
  output [3:0] io_in_0_b_bits_mask,
  output [31:0] io_in_0_b_bits_data,
  output  io_in_0_c_ready,
  input   io_in_0_c_valid,
  input  [2:0] io_in_0_c_bits_opcode,
  input  [2:0] io_in_0_c_bits_param,
  input  [2:0] io_in_0_c_bits_size,
  input  [4:0] io_in_0_c_bits_source,
  input  [28:0] io_in_0_c_bits_address,
  input  [31:0] io_in_0_c_bits_data,
  input   io_in_0_c_bits_error,
  input   io_in_0_d_ready,
  output  io_in_0_d_valid,
  output [2:0] io_in_0_d_bits_opcode,
  output [1:0] io_in_0_d_bits_param,
  output [2:0] io_in_0_d_bits_size,
  output [4:0] io_in_0_d_bits_source,
  output  io_in_0_d_bits_sink,
  output [1:0] io_in_0_d_bits_addr_lo,
  output [31:0] io_in_0_d_bits_data,
  output  io_in_0_d_bits_error,
  output  io_in_0_e_ready,
  input   io_in_0_e_valid,
  input   io_in_0_e_bits_sink,
  output  io_moff_hfclkrst,
  output  io_moff_corerst,
  output  io_wdog_rst,
  output  io_lfclk,
  output  io_pmu_vddpaden,
  output  io_pmu_padrst,
  input   io_pmu_dwakeup,
  input   io_lfextclk,
  input   io_resetCauses_wdogrst,
  input   io_resetCauses_erst,
  input   io_resetCauses_porrst
);
  wire  rtc_clock;
  wire  rtc_reset;
  wire  rtc_io_regs_cfg_write_valid;
  wire [31:0] rtc_io_regs_cfg_write_bits;
  wire [31:0] rtc_io_regs_cfg_read;
  wire  rtc_io_regs_countLo_write_valid;
  wire [31:0] rtc_io_regs_countLo_write_bits;
  wire [31:0] rtc_io_regs_countLo_read;
  wire  rtc_io_regs_countHi_write_valid;
  wire [31:0] rtc_io_regs_countHi_write_bits;
  wire [31:0] rtc_io_regs_countHi_read;
  wire  rtc_io_regs_s_write_valid;
  wire [31:0] rtc_io_regs_s_write_bits;
  wire [31:0] rtc_io_regs_s_read;
  wire  rtc_io_regs_cmp_0_write_valid;
  wire [31:0] rtc_io_regs_cmp_0_write_bits;
  wire [31:0] rtc_io_regs_cmp_0_read;
  wire  rtc_io_regs_feed_write_valid;
  wire [31:0] rtc_io_regs_feed_write_bits;
  wire [31:0] rtc_io_regs_feed_read;
  wire  rtc_io_regs_key_write_valid;
  wire [31:0] rtc_io_regs_key_write_bits;
  wire [31:0] rtc_io_regs_key_read;
  wire  rtc_io_ip_0;
  wire  pmu_clock;
  wire  pmu_reset;
  wire  pmu_io_wakeup_awakeup;
  wire  pmu_io_wakeup_dwakeup;
  wire  pmu_io_wakeup_rtc;
  wire  pmu_io_wakeup_reset;
  wire  pmu_io_control_hfclkrst;
  wire  pmu_io_control_corerst;
  wire  pmu_io_control_reserved1;
  wire  pmu_io_control_vddpaden;
  wire  pmu_io_control_reserved0;
  wire  pmu_io_regs_ie_write_valid;
  wire [3:0] pmu_io_regs_ie_write_bits;
  wire [3:0] pmu_io_regs_ie_read;
  wire  pmu_io_regs_cause_write_valid;
  wire [31:0] pmu_io_regs_cause_write_bits;
  wire [31:0] pmu_io_regs_cause_read;
  wire  pmu_io_regs_sleep_write_valid;
  wire [31:0] pmu_io_regs_sleep_write_bits;
  wire [31:0] pmu_io_regs_sleep_read;
  wire  pmu_io_regs_key_write_valid;
  wire [31:0] pmu_io_regs_key_write_bits;
  wire [31:0] pmu_io_regs_key_read;
  wire  pmu_io_regs_wakeupProgram_0_write_valid;
  wire [31:0] pmu_io_regs_wakeupProgram_0_write_bits;
  wire [31:0] pmu_io_regs_wakeupProgram_0_read;
  wire  pmu_io_regs_wakeupProgram_1_write_valid;
  wire [31:0] pmu_io_regs_wakeupProgram_1_write_bits;
  wire [31:0] pmu_io_regs_wakeupProgram_1_read;
  wire  pmu_io_regs_wakeupProgram_2_write_valid;
  wire [31:0] pmu_io_regs_wakeupProgram_2_write_bits;
  wire [31:0] pmu_io_regs_wakeupProgram_2_read;
  wire  pmu_io_regs_wakeupProgram_3_write_valid;
  wire [31:0] pmu_io_regs_wakeupProgram_3_write_bits;
  wire [31:0] pmu_io_regs_wakeupProgram_3_read;
  wire  pmu_io_regs_wakeupProgram_4_write_valid;
  wire [31:0] pmu_io_regs_wakeupProgram_4_write_bits;
  wire [31:0] pmu_io_regs_wakeupProgram_4_read;
  wire  pmu_io_regs_wakeupProgram_5_write_valid;
  wire [31:0] pmu_io_regs_wakeupProgram_5_write_bits;
  wire [31:0] pmu_io_regs_wakeupProgram_5_read;
  wire  pmu_io_regs_wakeupProgram_6_write_valid;
  wire [31:0] pmu_io_regs_wakeupProgram_6_write_bits;
  wire [31:0] pmu_io_regs_wakeupProgram_6_read;
  wire  pmu_io_regs_wakeupProgram_7_write_valid;
  wire [31:0] pmu_io_regs_wakeupProgram_7_write_bits;
  wire [31:0] pmu_io_regs_wakeupProgram_7_read;
  wire  pmu_io_regs_sleepProgram_0_write_valid;
  wire [31:0] pmu_io_regs_sleepProgram_0_write_bits;
  wire [31:0] pmu_io_regs_sleepProgram_0_read;
  wire  pmu_io_regs_sleepProgram_1_write_valid;
  wire [31:0] pmu_io_regs_sleepProgram_1_write_bits;
  wire [31:0] pmu_io_regs_sleepProgram_1_read;
  wire  pmu_io_regs_sleepProgram_2_write_valid;
  wire [31:0] pmu_io_regs_sleepProgram_2_write_bits;
  wire [31:0] pmu_io_regs_sleepProgram_2_read;
  wire  pmu_io_regs_sleepProgram_3_write_valid;
  wire [31:0] pmu_io_regs_sleepProgram_3_write_bits;
  wire [31:0] pmu_io_regs_sleepProgram_3_read;
  wire  pmu_io_regs_sleepProgram_4_write_valid;
  wire [31:0] pmu_io_regs_sleepProgram_4_write_bits;
  wire [31:0] pmu_io_regs_sleepProgram_4_read;
  wire  pmu_io_regs_sleepProgram_5_write_valid;
  wire [31:0] pmu_io_regs_sleepProgram_5_write_bits;
  wire [31:0] pmu_io_regs_sleepProgram_5_read;
  wire  pmu_io_regs_sleepProgram_6_write_valid;
  wire [31:0] pmu_io_regs_sleepProgram_6_write_bits;
  wire [31:0] pmu_io_regs_sleepProgram_6_read;
  wire  pmu_io_regs_sleepProgram_7_write_valid;
  wire [31:0] pmu_io_regs_sleepProgram_7_write_bits;
  wire [31:0] pmu_io_regs_sleepProgram_7_read;
  wire  pmu_io_resetCauses_wdogrst;
  wire  pmu_io_resetCauses_erst;
  wire  pmu_io_resetCauses_porrst;
  wire  wdog_clock;
  wire  wdog_reset;
  wire  wdog_io_regs_cfg_write_valid;
  wire [31:0] wdog_io_regs_cfg_write_bits;
  wire [31:0] wdog_io_regs_cfg_read;
  wire  wdog_io_regs_countLo_write_valid;
  wire [31:0] wdog_io_regs_countLo_write_bits;
  wire [31:0] wdog_io_regs_countLo_read;
  wire  wdog_io_regs_countHi_write_valid;
  wire [31:0] wdog_io_regs_countHi_write_bits;
  wire [31:0] wdog_io_regs_countHi_read;
  wire  wdog_io_regs_s_write_valid;
  wire [15:0] wdog_io_regs_s_write_bits;
  wire [15:0] wdog_io_regs_s_read;
  wire  wdog_io_regs_cmp_0_write_valid;
  wire [15:0] wdog_io_regs_cmp_0_write_bits;
  wire [15:0] wdog_io_regs_cmp_0_read;
  wire  wdog_io_regs_feed_write_valid;
  wire [31:0] wdog_io_regs_feed_write_bits;
  wire [31:0] wdog_io_regs_feed_read;
  wire  wdog_io_regs_key_write_valid;
  wire [31:0] wdog_io_regs_key_write_bits;
  wire [31:0] wdog_io_regs_key_read;
  wire  wdog_io_ip_0;
  wire  wdog_io_corerst;
  wire  wdog_io_rst;
  reg [31:0] backupRegs_0;
  reg [31:0] GEN_792;
  reg [31:0] backupRegs_1;
  reg [31:0] GEN_793;
  reg [31:0] backupRegs_2;
  reg [31:0] GEN_794;
  reg [31:0] backupRegs_3;
  reg [31:0] GEN_795;
  reg [31:0] backupRegs_4;
  reg [31:0] GEN_796;
  reg [31:0] backupRegs_5;
  reg [31:0] GEN_797;
  reg [31:0] backupRegs_6;
  reg [31:0] GEN_798;
  reg [31:0] backupRegs_7;
  reg [31:0] GEN_799;
  reg [31:0] backupRegs_8;
  reg [31:0] GEN_800;
  reg [31:0] backupRegs_9;
  reg [31:0] GEN_801;
  reg [31:0] backupRegs_10;
  reg [31:0] GEN_802;
  reg [31:0] backupRegs_11;
  reg [31:0] GEN_803;
  reg [31:0] backupRegs_12;
  reg [31:0] GEN_804;
  reg [31:0] backupRegs_13;
  reg [31:0] GEN_805;
  reg [31:0] backupRegs_14;
  reg [31:0] GEN_806;
  reg [31:0] backupRegs_15;
  reg [31:0] GEN_807;
  wire  T_953_ready;
  wire  T_953_valid;
  wire  T_953_bits_read;
  wire [9:0] T_953_bits_index;
  wire [31:0] T_953_bits_data;
  wire [3:0] T_953_bits_mask;
  wire [9:0] T_953_bits_extra;
  wire  T_970;
  wire [26:0] T_971;
  wire [1:0] T_972;
  wire [6:0] T_973;
  wire [9:0] T_974;
  wire  T_992_ready;
  wire  T_992_valid;
  wire  T_992_bits_read;
  wire [31:0] T_992_bits_data;
  wire [9:0] T_992_bits_extra;
  wire  T_1028_ready;
  wire  T_1028_valid;
  wire  T_1028_bits_read;
  wire [9:0] T_1028_bits_index;
  wire [31:0] T_1028_bits_data;
  wire [3:0] T_1028_bits_mask;
  wire [9:0] T_1028_bits_extra;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire  Queue_1_io_enq_bits_read;
  wire [9:0] Queue_1_io_enq_bits_index;
  wire [31:0] Queue_1_io_enq_bits_data;
  wire [3:0] Queue_1_io_enq_bits_mask;
  wire [9:0] Queue_1_io_enq_bits_extra;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire  Queue_1_io_deq_bits_read;
  wire [9:0] Queue_1_io_deq_bits_index;
  wire [31:0] Queue_1_io_deq_bits_data;
  wire [3:0] Queue_1_io_deq_bits_mask;
  wire [9:0] Queue_1_io_deq_bits_extra;
  wire  Queue_1_io_count;
  wire [9:0] T_1310;
  wire [9:0] T_1311;
  wire  T_1313;
  wire [9:0] T_1314;
  wire [9:0] T_1315;
  wire  T_1317;
  wire [9:0] T_1320;
  wire  T_1322;
  wire [9:0] T_1323;
  wire [9:0] T_1324;
  wire  T_1326;
  wire [9:0] T_1328;
  wire [9:0] T_1329;
  wire  T_1331;
  wire [9:0] T_1332;
  wire [9:0] T_1333;
  wire  T_1335;
  wire [9:0] T_1337;
  wire [9:0] T_1338;
  wire  T_1340;
  wire [9:0] T_1341;
  wire [9:0] T_1342;
  wire  T_1344;
  wire [9:0] T_1346;
  wire [9:0] T_1347;
  wire  T_1349;
  wire [9:0] T_1350;
  wire [9:0] T_1351;
  wire  T_1353;
  wire [9:0] T_1355;
  wire [9:0] T_1356;
  wire  T_1358;
  wire [9:0] T_1359;
  wire [9:0] T_1360;
  wire  T_1362;
  wire [9:0] T_1364;
  wire [9:0] T_1365;
  wire  T_1367;
  wire [9:0] T_1368;
  wire [9:0] T_1369;
  wire  T_1371;
  wire [9:0] T_1373;
  wire [9:0] T_1374;
  wire  T_1376;
  wire [9:0] T_1377;
  wire [9:0] T_1378;
  wire  T_1380;
  wire [9:0] T_1382;
  wire [9:0] T_1383;
  wire  T_1385;
  wire [9:0] T_1386;
  wire [9:0] T_1387;
  wire  T_1389;
  wire [9:0] T_1391;
  wire [9:0] T_1392;
  wire  T_1394;
  wire [9:0] T_1395;
  wire [9:0] T_1396;
  wire  T_1398;
  wire [9:0] T_1400;
  wire [9:0] T_1401;
  wire  T_1403;
  wire [9:0] T_1404;
  wire [9:0] T_1405;
  wire  T_1407;
  wire [9:0] T_1409;
  wire [9:0] T_1410;
  wire  T_1412;
  wire [9:0] T_1413;
  wire [9:0] T_1414;
  wire  T_1416;
  wire [9:0] T_1418;
  wire [9:0] T_1419;
  wire  T_1421;
  wire [9:0] T_1422;
  wire [9:0] T_1423;
  wire  T_1425;
  wire [9:0] T_1427;
  wire [9:0] T_1428;
  wire  T_1430;
  wire [9:0] T_1431;
  wire [9:0] T_1432;
  wire  T_1434;
  wire [9:0] T_1436;
  wire [9:0] T_1437;
  wire  T_1439;
  wire [9:0] T_1440;
  wire [9:0] T_1441;
  wire  T_1443;
  wire [9:0] T_1445;
  wire [9:0] T_1446;
  wire  T_1448;
  wire [9:0] T_1449;
  wire [9:0] T_1450;
  wire  T_1452;
  wire [9:0] T_1454;
  wire [9:0] T_1455;
  wire  T_1457;
  wire [9:0] T_1458;
  wire [9:0] T_1459;
  wire  T_1461;
  wire [9:0] T_1463;
  wire [9:0] T_1464;
  wire  T_1466;
  wire [9:0] T_1467;
  wire [9:0] T_1468;
  wire  T_1470;
  wire [9:0] T_1472;
  wire [9:0] T_1473;
  wire  T_1475;
  wire [9:0] T_1476;
  wire [9:0] T_1477;
  wire  T_1479;
  wire [9:0] T_1481;
  wire [9:0] T_1482;
  wire  T_1484;
  wire [9:0] T_1485;
  wire [9:0] T_1486;
  wire  T_1488;
  wire [9:0] T_1490;
  wire [9:0] T_1491;
  wire  T_1493;
  wire [9:0] T_1494;
  wire [9:0] T_1495;
  wire  T_1497;
  wire [9:0] T_1499;
  wire [9:0] T_1500;
  wire  T_1502;
  wire [9:0] T_1503;
  wire [9:0] T_1504;
  wire  T_1506;
  wire [9:0] T_1508;
  wire [9:0] T_1509;
  wire  T_1511;
  wire [9:0] T_1512;
  wire [9:0] T_1513;
  wire  T_1515;
  wire [9:0] T_1517;
  wire [9:0] T_1518;
  wire  T_1520;
  wire [9:0] T_1521;
  wire [9:0] T_1522;
  wire  T_1524;
  wire [9:0] T_1526;
  wire [9:0] T_1527;
  wire  T_1529;
  wire [9:0] T_1530;
  wire [9:0] T_1531;
  wire  T_1533;
  wire [9:0] T_1535;
  wire [9:0] T_1536;
  wire  T_1538;
  wire [9:0] T_1539;
  wire [9:0] T_1540;
  wire  T_1542;
  wire [9:0] T_1544;
  wire [9:0] T_1545;
  wire  T_1547;
  wire [9:0] T_1548;
  wire [9:0] T_1549;
  wire  T_1551;
  wire [9:0] T_1553;
  wire [9:0] T_1554;
  wire  T_1556;
  wire [9:0] T_1557;
  wire [9:0] T_1558;
  wire  T_1560;
  wire [9:0] T_1562;
  wire [9:0] T_1563;
  wire  T_1565;
  wire [9:0] T_1566;
  wire [9:0] T_1567;
  wire  T_1569;
  wire [9:0] T_1571;
  wire [9:0] T_1572;
  wire  T_1574;
  wire [9:0] T_1575;
  wire [9:0] T_1576;
  wire  T_1578;
  wire [9:0] T_1580;
  wire [9:0] T_1581;
  wire  T_1583;
  wire [9:0] T_1584;
  wire [9:0] T_1585;
  wire  T_1587;
  wire [9:0] T_1589;
  wire [9:0] T_1590;
  wire  T_1592;
  wire [9:0] T_1593;
  wire [9:0] T_1594;
  wire  T_1596;
  wire [9:0] T_1598;
  wire [9:0] T_1599;
  wire  T_1601;
  wire [9:0] T_1602;
  wire [9:0] T_1603;
  wire  T_1605;
  wire [9:0] T_1607;
  wire [9:0] T_1608;
  wire  T_1610;
  wire [9:0] T_1611;
  wire [9:0] T_1612;
  wire  T_1614;
  wire [9:0] T_1616;
  wire [9:0] T_1617;
  wire  T_1619;
  wire [9:0] T_1620;
  wire [9:0] T_1621;
  wire  T_1623;
  wire [9:0] T_1625;
  wire [9:0] T_1626;
  wire  T_1628;
  wire [9:0] T_1629;
  wire [9:0] T_1630;
  wire  T_1632;
  wire [9:0] T_1634;
  wire [9:0] T_1635;
  wire  T_1637;
  wire [9:0] T_1638;
  wire [9:0] T_1639;
  wire  T_1641;
  wire [9:0] T_1643;
  wire [9:0] T_1644;
  wire  T_1646;
  wire [9:0] T_1647;
  wire [9:0] T_1648;
  wire  T_1650;
  wire [9:0] T_1652;
  wire [9:0] T_1653;
  wire  T_1655;
  wire [9:0] T_1656;
  wire [9:0] T_1657;
  wire  T_1659;
  wire [9:0] T_1661;
  wire [9:0] T_1662;
  wire  T_1664;
  wire [9:0] T_1665;
  wire [9:0] T_1666;
  wire  T_1668;
  wire [9:0] T_1670;
  wire [9:0] T_1671;
  wire  T_1673;
  wire [9:0] T_1674;
  wire [9:0] T_1675;
  wire  T_1677;
  wire [9:0] T_1679;
  wire [9:0] T_1680;
  wire  T_1682;
  wire [9:0] T_1683;
  wire [9:0] T_1684;
  wire  T_1686;
  wire [9:0] T_1688;
  wire [9:0] T_1689;
  wire  T_1691;
  wire [9:0] T_1692;
  wire [9:0] T_1693;
  wire  T_1695;
  wire [9:0] T_1697;
  wire [9:0] T_1698;
  wire  T_1700;
  wire [9:0] T_1701;
  wire [9:0] T_1702;
  wire  T_1704;
  wire [9:0] T_1706;
  wire [9:0] T_1707;
  wire  T_1709;
  wire [9:0] T_1710;
  wire [9:0] T_1711;
  wire  T_1713;
  wire [9:0] T_1715;
  wire [9:0] T_1716;
  wire  T_1718;
  wire [9:0] T_1719;
  wire [9:0] T_1720;
  wire  T_1722;
  wire [9:0] T_1724;
  wire [9:0] T_1725;
  wire  T_1727;
  wire [9:0] T_1728;
  wire [9:0] T_1729;
  wire  T_1731;
  wire [9:0] T_1733;
  wire [9:0] T_1734;
  wire  T_1736;
  wire [9:0] T_1737;
  wire [9:0] T_1738;
  wire  T_1740;
  wire [9:0] T_1742;
  wire [9:0] T_1743;
  wire  T_1745;
  wire [9:0] T_1746;
  wire [9:0] T_1747;
  wire  T_1749;
  wire [9:0] T_1751;
  wire [9:0] T_1752;
  wire  T_1754;
  wire [9:0] T_1755;
  wire [9:0] T_1756;
  wire  T_1758;
  wire  T_1762_0;
  wire  T_1762_1;
  wire  T_1762_2;
  wire  T_1762_3;
  wire  T_1762_4;
  wire  T_1762_5;
  wire  T_1762_6;
  wire  T_1762_7;
  wire  T_1762_8;
  wire  T_1762_9;
  wire  T_1762_10;
  wire  T_1762_11;
  wire  T_1762_12;
  wire  T_1762_13;
  wire  T_1762_14;
  wire  T_1762_15;
  wire  T_1762_16;
  wire  T_1762_17;
  wire  T_1762_18;
  wire  T_1762_19;
  wire  T_1762_20;
  wire  T_1762_21;
  wire  T_1762_22;
  wire  T_1762_23;
  wire  T_1762_24;
  wire  T_1762_25;
  wire  T_1762_26;
  wire  T_1762_27;
  wire  T_1762_28;
  wire  T_1762_29;
  wire  T_1762_30;
  wire  T_1762_31;
  wire  T_1762_32;
  wire  T_1762_33;
  wire  T_1762_34;
  wire  T_1762_35;
  wire  T_1762_36;
  wire  T_1762_37;
  wire  T_1762_38;
  wire  T_1762_39;
  wire  T_1762_40;
  wire  T_1762_41;
  wire  T_1762_42;
  wire  T_1762_43;
  wire  T_1762_44;
  wire  T_1762_45;
  wire  T_1762_46;
  wire  T_1762_47;
  wire  T_1762_48;
  wire  T_1762_49;
  wire  T_1767_0;
  wire  T_1767_1;
  wire  T_1767_2;
  wire  T_1767_3;
  wire  T_1767_4;
  wire  T_1767_5;
  wire  T_1767_6;
  wire  T_1767_7;
  wire  T_1767_8;
  wire  T_1767_9;
  wire  T_1767_10;
  wire  T_1767_11;
  wire  T_1767_12;
  wire  T_1767_13;
  wire  T_1767_14;
  wire  T_1767_15;
  wire  T_1767_16;
  wire  T_1767_17;
  wire  T_1767_18;
  wire  T_1767_19;
  wire  T_1767_20;
  wire  T_1767_21;
  wire  T_1767_22;
  wire  T_1767_23;
  wire  T_1767_24;
  wire  T_1767_25;
  wire  T_1767_26;
  wire  T_1767_27;
  wire  T_1767_28;
  wire  T_1767_29;
  wire  T_1767_30;
  wire  T_1767_31;
  wire  T_1767_32;
  wire  T_1767_33;
  wire  T_1767_34;
  wire  T_1767_35;
  wire  T_1767_36;
  wire  T_1767_37;
  wire  T_1767_38;
  wire  T_1767_39;
  wire  T_1767_40;
  wire  T_1767_41;
  wire  T_1767_42;
  wire  T_1767_43;
  wire  T_1767_44;
  wire  T_1767_45;
  wire  T_1767_46;
  wire  T_1767_47;
  wire  T_1767_48;
  wire  T_1767_49;
  wire  T_1772_0;
  wire  T_1772_1;
  wire  T_1772_2;
  wire  T_1772_3;
  wire  T_1772_4;
  wire  T_1772_5;
  wire  T_1772_6;
  wire  T_1772_7;
  wire  T_1772_8;
  wire  T_1772_9;
  wire  T_1772_10;
  wire  T_1772_11;
  wire  T_1772_12;
  wire  T_1772_13;
  wire  T_1772_14;
  wire  T_1772_15;
  wire  T_1772_16;
  wire  T_1772_17;
  wire  T_1772_18;
  wire  T_1772_19;
  wire  T_1772_20;
  wire  T_1772_21;
  wire  T_1772_22;
  wire  T_1772_23;
  wire  T_1772_24;
  wire  T_1772_25;
  wire  T_1772_26;
  wire  T_1772_27;
  wire  T_1772_28;
  wire  T_1772_29;
  wire  T_1772_30;
  wire  T_1772_31;
  wire  T_1772_32;
  wire  T_1772_33;
  wire  T_1772_34;
  wire  T_1772_35;
  wire  T_1772_36;
  wire  T_1772_37;
  wire  T_1772_38;
  wire  T_1772_39;
  wire  T_1772_40;
  wire  T_1772_41;
  wire  T_1772_42;
  wire  T_1772_43;
  wire  T_1772_44;
  wire  T_1772_45;
  wire  T_1772_46;
  wire  T_1772_47;
  wire  T_1772_48;
  wire  T_1772_49;
  wire  T_1777_0;
  wire  T_1777_1;
  wire  T_1777_2;
  wire  T_1777_3;
  wire  T_1777_4;
  wire  T_1777_5;
  wire  T_1777_6;
  wire  T_1777_7;
  wire  T_1777_8;
  wire  T_1777_9;
  wire  T_1777_10;
  wire  T_1777_11;
  wire  T_1777_12;
  wire  T_1777_13;
  wire  T_1777_14;
  wire  T_1777_15;
  wire  T_1777_16;
  wire  T_1777_17;
  wire  T_1777_18;
  wire  T_1777_19;
  wire  T_1777_20;
  wire  T_1777_21;
  wire  T_1777_22;
  wire  T_1777_23;
  wire  T_1777_24;
  wire  T_1777_25;
  wire  T_1777_26;
  wire  T_1777_27;
  wire  T_1777_28;
  wire  T_1777_29;
  wire  T_1777_30;
  wire  T_1777_31;
  wire  T_1777_32;
  wire  T_1777_33;
  wire  T_1777_34;
  wire  T_1777_35;
  wire  T_1777_36;
  wire  T_1777_37;
  wire  T_1777_38;
  wire  T_1777_39;
  wire  T_1777_40;
  wire  T_1777_41;
  wire  T_1777_42;
  wire  T_1777_43;
  wire  T_1777_44;
  wire  T_1777_45;
  wire  T_1777_46;
  wire  T_1777_47;
  wire  T_1777_48;
  wire  T_1777_49;
  wire  T_1782_0;
  wire  T_1782_1;
  wire  T_1782_2;
  wire  T_1782_3;
  wire  T_1782_4;
  wire  T_1782_5;
  wire  T_1782_6;
  wire  T_1782_7;
  wire  T_1782_8;
  wire  T_1782_9;
  wire  T_1782_10;
  wire  T_1782_11;
  wire  T_1782_12;
  wire  T_1782_13;
  wire  T_1782_14;
  wire  T_1782_15;
  wire  T_1782_16;
  wire  T_1782_17;
  wire  T_1782_18;
  wire  T_1782_19;
  wire  T_1782_20;
  wire  T_1782_21;
  wire  T_1782_22;
  wire  T_1782_23;
  wire  T_1782_24;
  wire  T_1782_25;
  wire  T_1782_26;
  wire  T_1782_27;
  wire  T_1782_28;
  wire  T_1782_29;
  wire  T_1782_30;
  wire  T_1782_31;
  wire  T_1782_32;
  wire  T_1782_33;
  wire  T_1782_34;
  wire  T_1782_35;
  wire  T_1782_36;
  wire  T_1782_37;
  wire  T_1782_38;
  wire  T_1782_39;
  wire  T_1782_40;
  wire  T_1782_41;
  wire  T_1782_42;
  wire  T_1782_43;
  wire  T_1782_44;
  wire  T_1782_45;
  wire  T_1782_46;
  wire  T_1782_47;
  wire  T_1782_48;
  wire  T_1782_49;
  wire  T_1787_0;
  wire  T_1787_1;
  wire  T_1787_2;
  wire  T_1787_3;
  wire  T_1787_4;
  wire  T_1787_5;
  wire  T_1787_6;
  wire  T_1787_7;
  wire  T_1787_8;
  wire  T_1787_9;
  wire  T_1787_10;
  wire  T_1787_11;
  wire  T_1787_12;
  wire  T_1787_13;
  wire  T_1787_14;
  wire  T_1787_15;
  wire  T_1787_16;
  wire  T_1787_17;
  wire  T_1787_18;
  wire  T_1787_19;
  wire  T_1787_20;
  wire  T_1787_21;
  wire  T_1787_22;
  wire  T_1787_23;
  wire  T_1787_24;
  wire  T_1787_25;
  wire  T_1787_26;
  wire  T_1787_27;
  wire  T_1787_28;
  wire  T_1787_29;
  wire  T_1787_30;
  wire  T_1787_31;
  wire  T_1787_32;
  wire  T_1787_33;
  wire  T_1787_34;
  wire  T_1787_35;
  wire  T_1787_36;
  wire  T_1787_37;
  wire  T_1787_38;
  wire  T_1787_39;
  wire  T_1787_40;
  wire  T_1787_41;
  wire  T_1787_42;
  wire  T_1787_43;
  wire  T_1787_44;
  wire  T_1787_45;
  wire  T_1787_46;
  wire  T_1787_47;
  wire  T_1787_48;
  wire  T_1787_49;
  wire  T_1792_0;
  wire  T_1792_1;
  wire  T_1792_2;
  wire  T_1792_3;
  wire  T_1792_4;
  wire  T_1792_5;
  wire  T_1792_6;
  wire  T_1792_7;
  wire  T_1792_8;
  wire  T_1792_9;
  wire  T_1792_10;
  wire  T_1792_11;
  wire  T_1792_12;
  wire  T_1792_13;
  wire  T_1792_14;
  wire  T_1792_15;
  wire  T_1792_16;
  wire  T_1792_17;
  wire  T_1792_18;
  wire  T_1792_19;
  wire  T_1792_20;
  wire  T_1792_21;
  wire  T_1792_22;
  wire  T_1792_23;
  wire  T_1792_24;
  wire  T_1792_25;
  wire  T_1792_26;
  wire  T_1792_27;
  wire  T_1792_28;
  wire  T_1792_29;
  wire  T_1792_30;
  wire  T_1792_31;
  wire  T_1792_32;
  wire  T_1792_33;
  wire  T_1792_34;
  wire  T_1792_35;
  wire  T_1792_36;
  wire  T_1792_37;
  wire  T_1792_38;
  wire  T_1792_39;
  wire  T_1792_40;
  wire  T_1792_41;
  wire  T_1792_42;
  wire  T_1792_43;
  wire  T_1792_44;
  wire  T_1792_45;
  wire  T_1792_46;
  wire  T_1792_47;
  wire  T_1792_48;
  wire  T_1792_49;
  wire  T_1797_0;
  wire  T_1797_1;
  wire  T_1797_2;
  wire  T_1797_3;
  wire  T_1797_4;
  wire  T_1797_5;
  wire  T_1797_6;
  wire  T_1797_7;
  wire  T_1797_8;
  wire  T_1797_9;
  wire  T_1797_10;
  wire  T_1797_11;
  wire  T_1797_12;
  wire  T_1797_13;
  wire  T_1797_14;
  wire  T_1797_15;
  wire  T_1797_16;
  wire  T_1797_17;
  wire  T_1797_18;
  wire  T_1797_19;
  wire  T_1797_20;
  wire  T_1797_21;
  wire  T_1797_22;
  wire  T_1797_23;
  wire  T_1797_24;
  wire  T_1797_25;
  wire  T_1797_26;
  wire  T_1797_27;
  wire  T_1797_28;
  wire  T_1797_29;
  wire  T_1797_30;
  wire  T_1797_31;
  wire  T_1797_32;
  wire  T_1797_33;
  wire  T_1797_34;
  wire  T_1797_35;
  wire  T_1797_36;
  wire  T_1797_37;
  wire  T_1797_38;
  wire  T_1797_39;
  wire  T_1797_40;
  wire  T_1797_41;
  wire  T_1797_42;
  wire  T_1797_43;
  wire  T_1797_44;
  wire  T_1797_45;
  wire  T_1797_46;
  wire  T_1797_47;
  wire  T_1797_48;
  wire  T_1797_49;
  wire  T_2462;
  wire  T_2463;
  wire  T_2464;
  wire  T_2465;
  wire [7:0] T_2469;
  wire [7:0] T_2473;
  wire [7:0] T_2477;
  wire [7:0] T_2481;
  wire [15:0] T_2482;
  wire [15:0] T_2483;
  wire [31:0] T_2484;
  wire [31:0] T_2496;
  wire  T_2498;
  wire  T_2504;
  wire [31:0] T_2505;
  wire [31:0] T_2520;
  wire  T_2544;
  wire [31:0] T_2560;
  wire  T_2584;
  wire [31:0] GEN_6;
  wire  T_2624;
  wire [31:0] T_2640;
  wire  T_2664;
  wire [31:0] GEN_7;
  wire  T_2704;
  wire [31:0] T_2720;
  wire  T_2744;
  wire [31:0] GEN_8;
  wire  T_2784;
  wire [31:0] T_2800;
  wire  T_2824;
  wire [31:0] T_2840;
  wire  T_2864;
  wire [31:0] T_2880;
  wire  T_2904;
  wire [31:0] GEN_9;
  wire  T_2944;
  wire [31:0] T_2960;
  wire  T_2984;
  wire [31:0] GEN_10;
  wire  T_3024;
  wire [31:0] T_3040;
  wire  T_3064;
  wire [31:0] T_3080;
  wire  T_3104;
  wire [31:0] GEN_11;
  wire  T_3144;
  wire [31:0] T_3160;
  wire  T_3184;
  wire [31:0] T_3200;
  wire  T_3224;
  wire [31:0] GEN_12;
  wire  T_3264;
  wire [31:0] GEN_13;
  wire  T_3304;
  wire [31:0] GEN_14;
  wire  T_3344;
  wire [31:0] T_3360;
  wire  T_3384;
  wire [31:0] T_3400;
  wire  T_3424;
  wire [31:0] GEN_15;
  wire  T_3464;
  wire [31:0] T_3480;
  wire  T_3504;
  wire [31:0] T_3520;
  wire  T_3544;
  wire [31:0] T_3560;
  wire  T_3584;
  wire [31:0] T_3600;
  wire  T_3624;
  wire [31:0] GEN_16;
  wire  T_3664;
  wire [31:0] T_3680;
  wire  T_3704;
  wire [31:0] T_3720;
  wire [3:0] T_3732;
  wire [3:0] T_3736;
  wire  T_3738;
  wire  T_3744;
  wire [3:0] T_3745;
  wire [3:0] T_3760;
  wire  T_3784;
  wire [31:0] GEN_17;
  wire  T_3824;
  wire [31:0] T_3840;
  wire  T_3864;
  wire [31:0] T_3880;
  wire  T_3904;
  wire [31:0] T_3920;
  wire  T_3944;
  wire [31:0] T_3960;
  wire  T_3984;
  wire [31:0] GEN_18;
  wire  T_4024;
  wire [31:0] GEN_19;
  wire  T_4064;
  wire [31:0] T_4080;
  wire [15:0] T_4092;
  wire [15:0] T_4096;
  wire  T_4098;
  wire  T_4104;
  wire [15:0] T_4105;
  wire [15:0] T_4120;
  wire  T_4144;
  wire [31:0] T_4160;
  wire  T_4184;
  wire [31:0] T_4200;
  wire  T_4224;
  wire [31:0] GEN_20;
  wire  T_4264;
  wire [31:0] T_4280;
  wire  T_4304;
  wire [15:0] T_4320;
  wire  T_4344;
  wire [31:0] T_4360;
  wire  T_4384;
  wire [31:0] GEN_21;
  wire  T_4424;
  wire [31:0] T_4440;
  wire  T_4464;
  wire [31:0] T_4480;
  wire  T_4486;
  wire  T_4488;
  wire  T_4493;
  wire  T_4495;
  wire  T_4497;
  wire  T_4499;
  wire  T_4501;
  wire  T_4503;
  wire  T_4508;
  wire  T_4510;
  wire  T_4512;
  wire  T_4514;
  wire  T_4516;
  wire  T_4518;
  wire  T_4541;
  wire  T_4543;
  wire  T_4548;
  wire  T_4550;
  wire  T_4552;
  wire  T_4554;
  wire  T_4556;
  wire  T_4558;
  wire  T_4563;
  wire  T_4565;
  wire  T_4567;
  wire  T_4569;
  wire  T_4571;
  wire  T_4573;
  wire  T_4596;
  wire  T_4598;
  wire  T_4600;
  wire  T_4602;
  wire  T_4604;
  wire  T_4606;
  wire  T_4608;
  wire  T_4610;
  wire  T_4612;
  wire  T_4614;
  wire  T_4616;
  wire  T_4618;
  wire  T_4620;
  wire  T_4622;
  wire  T_4624;
  wire  T_4626;
  wire  T_4628;
  wire  T_4630;
  wire  T_4632;
  wire  T_4634;
  wire  T_4636;
  wire  T_4638;
  wire  T_4640;
  wire  T_4642;
  wire  T_4644;
  wire  T_4646;
  wire  T_4648;
  wire  T_4650;
  wire  T_4652;
  wire  T_4654;
  wire  T_4656;
  wire  T_4658;
  wire  T_4708;
  wire  T_4710;
  wire  T_4712;
  wire  T_4714;
  wire  T_4716;
  wire  T_4718;
  wire  T_4720;
  wire  T_4722;
  wire  T_4724;
  wire  T_4726;
  wire  T_4728;
  wire  T_4730;
  wire  T_4732;
  wire  T_4734;
  wire  T_4736;
  wire  T_4738;
  wire  T_4740;
  wire  T_4742;
  wire  T_4744;
  wire  T_4746;
  wire  T_4748;
  wire  T_4750;
  wire  T_4752;
  wire  T_4754;
  wire  T_4756;
  wire  T_4758;
  wire  T_4760;
  wire  T_4762;
  wire  T_4764;
  wire  T_4766;
  wire  T_4768;
  wire  T_4770;
  wire  T_4772;
  wire  T_4774;
  wire  T_4776;
  wire  T_4778;
  wire  T_4780;
  wire  T_4782;
  wire  T_4784;
  wire  T_4786;
  wire  T_5050_0;
  wire  T_5050_1;
  wire  T_5050_2;
  wire  T_5050_3;
  wire  T_5050_4;
  wire  T_5050_5;
  wire  T_5050_6;
  wire  T_5050_7;
  wire  T_5050_8;
  wire  T_5050_9;
  wire  T_5050_10;
  wire  T_5050_11;
  wire  T_5050_12;
  wire  T_5050_13;
  wire  T_5050_14;
  wire  T_5050_15;
  wire  T_5050_16;
  wire  T_5050_17;
  wire  T_5050_18;
  wire  T_5050_19;
  wire  T_5050_20;
  wire  T_5050_21;
  wire  T_5050_22;
  wire  T_5050_23;
  wire  T_5050_24;
  wire  T_5050_25;
  wire  T_5050_26;
  wire  T_5050_27;
  wire  T_5050_28;
  wire  T_5050_29;
  wire  T_5050_30;
  wire  T_5050_31;
  wire  T_5050_32;
  wire  T_5050_33;
  wire  T_5050_34;
  wire  T_5050_35;
  wire  T_5050_36;
  wire  T_5050_37;
  wire  T_5050_38;
  wire  T_5050_39;
  wire  T_5050_40;
  wire  T_5050_41;
  wire  T_5050_42;
  wire  T_5050_43;
  wire  T_5050_44;
  wire  T_5050_45;
  wire  T_5050_46;
  wire  T_5050_47;
  wire  T_5050_48;
  wire  T_5050_49;
  wire  T_5050_50;
  wire  T_5050_51;
  wire  T_5050_52;
  wire  T_5050_53;
  wire  T_5050_54;
  wire  T_5050_55;
  wire  T_5050_56;
  wire  T_5050_57;
  wire  T_5050_58;
  wire  T_5050_59;
  wire  T_5050_60;
  wire  T_5050_61;
  wire  T_5050_62;
  wire  T_5050_63;
  wire  T_5050_64;
  wire  T_5050_65;
  wire  T_5050_66;
  wire  T_5050_67;
  wire  T_5050_68;
  wire  T_5050_69;
  wire  T_5050_70;
  wire  T_5050_71;
  wire  T_5050_72;
  wire  T_5050_73;
  wire  T_5050_74;
  wire  T_5050_75;
  wire  T_5050_76;
  wire  T_5050_77;
  wire  T_5050_78;
  wire  T_5050_79;
  wire  T_5050_80;
  wire  T_5050_81;
  wire  T_5050_82;
  wire  T_5050_83;
  wire  T_5050_84;
  wire  T_5050_85;
  wire  T_5050_86;
  wire  T_5050_87;
  wire  T_5050_88;
  wire  T_5050_89;
  wire  T_5050_90;
  wire  T_5050_91;
  wire  T_5050_92;
  wire  T_5050_93;
  wire  T_5050_94;
  wire  T_5050_95;
  wire  T_5050_96;
  wire  T_5050_97;
  wire  T_5050_98;
  wire  T_5050_99;
  wire  T_5050_100;
  wire  T_5050_101;
  wire  T_5050_102;
  wire  T_5050_103;
  wire  T_5050_104;
  wire  T_5050_105;
  wire  T_5050_106;
  wire  T_5050_107;
  wire  T_5050_108;
  wire  T_5050_109;
  wire  T_5050_110;
  wire  T_5050_111;
  wire  T_5050_112;
  wire  T_5050_113;
  wire  T_5050_114;
  wire  T_5050_115;
  wire  T_5050_116;
  wire  T_5050_117;
  wire  T_5050_118;
  wire  T_5050_119;
  wire  T_5050_120;
  wire  T_5050_121;
  wire  T_5050_122;
  wire  T_5050_123;
  wire  T_5050_124;
  wire  T_5050_125;
  wire  T_5050_126;
  wire  T_5050_127;
  wire  T_5184;
  wire  T_5191;
  wire  T_5195;
  wire  T_5199;
  wire  T_5206;
  wire  T_5210;
  wire  T_5214;
  wire  T_5239;
  wire  T_5246;
  wire  T_5250;
  wire  T_5254;
  wire  T_5261;
  wire  T_5265;
  wire  T_5269;
  wire  T_5294;
  wire  T_5298;
  wire  T_5302;
  wire  T_5306;
  wire  T_5310;
  wire  T_5314;
  wire  T_5318;
  wire  T_5322;
  wire  T_5326;
  wire  T_5330;
  wire  T_5334;
  wire  T_5338;
  wire  T_5342;
  wire  T_5346;
  wire  T_5350;
  wire  T_5354;
  wire  T_5406;
  wire  T_5410;
  wire  T_5414;
  wire  T_5418;
  wire  T_5422;
  wire  T_5426;
  wire  T_5430;
  wire  T_5434;
  wire  T_5438;
  wire  T_5442;
  wire  T_5446;
  wire  T_5450;
  wire  T_5454;
  wire  T_5458;
  wire  T_5462;
  wire  T_5466;
  wire  T_5470;
  wire  T_5474;
  wire  T_5478;
  wire  T_5482;
  wire  T_5746_0;
  wire  T_5746_1;
  wire  T_5746_2;
  wire  T_5746_3;
  wire  T_5746_4;
  wire  T_5746_5;
  wire  T_5746_6;
  wire  T_5746_7;
  wire  T_5746_8;
  wire  T_5746_9;
  wire  T_5746_10;
  wire  T_5746_11;
  wire  T_5746_12;
  wire  T_5746_13;
  wire  T_5746_14;
  wire  T_5746_15;
  wire  T_5746_16;
  wire  T_5746_17;
  wire  T_5746_18;
  wire  T_5746_19;
  wire  T_5746_20;
  wire  T_5746_21;
  wire  T_5746_22;
  wire  T_5746_23;
  wire  T_5746_24;
  wire  T_5746_25;
  wire  T_5746_26;
  wire  T_5746_27;
  wire  T_5746_28;
  wire  T_5746_29;
  wire  T_5746_30;
  wire  T_5746_31;
  wire  T_5746_32;
  wire  T_5746_33;
  wire  T_5746_34;
  wire  T_5746_35;
  wire  T_5746_36;
  wire  T_5746_37;
  wire  T_5746_38;
  wire  T_5746_39;
  wire  T_5746_40;
  wire  T_5746_41;
  wire  T_5746_42;
  wire  T_5746_43;
  wire  T_5746_44;
  wire  T_5746_45;
  wire  T_5746_46;
  wire  T_5746_47;
  wire  T_5746_48;
  wire  T_5746_49;
  wire  T_5746_50;
  wire  T_5746_51;
  wire  T_5746_52;
  wire  T_5746_53;
  wire  T_5746_54;
  wire  T_5746_55;
  wire  T_5746_56;
  wire  T_5746_57;
  wire  T_5746_58;
  wire  T_5746_59;
  wire  T_5746_60;
  wire  T_5746_61;
  wire  T_5746_62;
  wire  T_5746_63;
  wire  T_5746_64;
  wire  T_5746_65;
  wire  T_5746_66;
  wire  T_5746_67;
  wire  T_5746_68;
  wire  T_5746_69;
  wire  T_5746_70;
  wire  T_5746_71;
  wire  T_5746_72;
  wire  T_5746_73;
  wire  T_5746_74;
  wire  T_5746_75;
  wire  T_5746_76;
  wire  T_5746_77;
  wire  T_5746_78;
  wire  T_5746_79;
  wire  T_5746_80;
  wire  T_5746_81;
  wire  T_5746_82;
  wire  T_5746_83;
  wire  T_5746_84;
  wire  T_5746_85;
  wire  T_5746_86;
  wire  T_5746_87;
  wire  T_5746_88;
  wire  T_5746_89;
  wire  T_5746_90;
  wire  T_5746_91;
  wire  T_5746_92;
  wire  T_5746_93;
  wire  T_5746_94;
  wire  T_5746_95;
  wire  T_5746_96;
  wire  T_5746_97;
  wire  T_5746_98;
  wire  T_5746_99;
  wire  T_5746_100;
  wire  T_5746_101;
  wire  T_5746_102;
  wire  T_5746_103;
  wire  T_5746_104;
  wire  T_5746_105;
  wire  T_5746_106;
  wire  T_5746_107;
  wire  T_5746_108;
  wire  T_5746_109;
  wire  T_5746_110;
  wire  T_5746_111;
  wire  T_5746_112;
  wire  T_5746_113;
  wire  T_5746_114;
  wire  T_5746_115;
  wire  T_5746_116;
  wire  T_5746_117;
  wire  T_5746_118;
  wire  T_5746_119;
  wire  T_5746_120;
  wire  T_5746_121;
  wire  T_5746_122;
  wire  T_5746_123;
  wire  T_5746_124;
  wire  T_5746_125;
  wire  T_5746_126;
  wire  T_5746_127;
  wire  T_5878;
  wire  T_5880;
  wire  T_5885;
  wire  T_5887;
  wire  T_5889;
  wire  T_5891;
  wire  T_5893;
  wire  T_5895;
  wire  T_5900;
  wire  T_5902;
  wire  T_5904;
  wire  T_5906;
  wire  T_5908;
  wire  T_5910;
  wire  T_5933;
  wire  T_5935;
  wire  T_5940;
  wire  T_5942;
  wire  T_5944;
  wire  T_5946;
  wire  T_5948;
  wire  T_5950;
  wire  T_5955;
  wire  T_5957;
  wire  T_5959;
  wire  T_5961;
  wire  T_5963;
  wire  T_5965;
  wire  T_5988;
  wire  T_5990;
  wire  T_5992;
  wire  T_5994;
  wire  T_5996;
  wire  T_5998;
  wire  T_6000;
  wire  T_6002;
  wire  T_6004;
  wire  T_6006;
  wire  T_6008;
  wire  T_6010;
  wire  T_6012;
  wire  T_6014;
  wire  T_6016;
  wire  T_6018;
  wire  T_6020;
  wire  T_6022;
  wire  T_6024;
  wire  T_6026;
  wire  T_6028;
  wire  T_6030;
  wire  T_6032;
  wire  T_6034;
  wire  T_6036;
  wire  T_6038;
  wire  T_6040;
  wire  T_6042;
  wire  T_6044;
  wire  T_6046;
  wire  T_6048;
  wire  T_6050;
  wire  T_6100;
  wire  T_6102;
  wire  T_6104;
  wire  T_6106;
  wire  T_6108;
  wire  T_6110;
  wire  T_6112;
  wire  T_6114;
  wire  T_6116;
  wire  T_6118;
  wire  T_6120;
  wire  T_6122;
  wire  T_6124;
  wire  T_6126;
  wire  T_6128;
  wire  T_6130;
  wire  T_6132;
  wire  T_6134;
  wire  T_6136;
  wire  T_6138;
  wire  T_6140;
  wire  T_6142;
  wire  T_6144;
  wire  T_6146;
  wire  T_6148;
  wire  T_6150;
  wire  T_6152;
  wire  T_6154;
  wire  T_6156;
  wire  T_6158;
  wire  T_6160;
  wire  T_6162;
  wire  T_6164;
  wire  T_6166;
  wire  T_6168;
  wire  T_6170;
  wire  T_6172;
  wire  T_6174;
  wire  T_6176;
  wire  T_6178;
  wire  T_6442_0;
  wire  T_6442_1;
  wire  T_6442_2;
  wire  T_6442_3;
  wire  T_6442_4;
  wire  T_6442_5;
  wire  T_6442_6;
  wire  T_6442_7;
  wire  T_6442_8;
  wire  T_6442_9;
  wire  T_6442_10;
  wire  T_6442_11;
  wire  T_6442_12;
  wire  T_6442_13;
  wire  T_6442_14;
  wire  T_6442_15;
  wire  T_6442_16;
  wire  T_6442_17;
  wire  T_6442_18;
  wire  T_6442_19;
  wire  T_6442_20;
  wire  T_6442_21;
  wire  T_6442_22;
  wire  T_6442_23;
  wire  T_6442_24;
  wire  T_6442_25;
  wire  T_6442_26;
  wire  T_6442_27;
  wire  T_6442_28;
  wire  T_6442_29;
  wire  T_6442_30;
  wire  T_6442_31;
  wire  T_6442_32;
  wire  T_6442_33;
  wire  T_6442_34;
  wire  T_6442_35;
  wire  T_6442_36;
  wire  T_6442_37;
  wire  T_6442_38;
  wire  T_6442_39;
  wire  T_6442_40;
  wire  T_6442_41;
  wire  T_6442_42;
  wire  T_6442_43;
  wire  T_6442_44;
  wire  T_6442_45;
  wire  T_6442_46;
  wire  T_6442_47;
  wire  T_6442_48;
  wire  T_6442_49;
  wire  T_6442_50;
  wire  T_6442_51;
  wire  T_6442_52;
  wire  T_6442_53;
  wire  T_6442_54;
  wire  T_6442_55;
  wire  T_6442_56;
  wire  T_6442_57;
  wire  T_6442_58;
  wire  T_6442_59;
  wire  T_6442_60;
  wire  T_6442_61;
  wire  T_6442_62;
  wire  T_6442_63;
  wire  T_6442_64;
  wire  T_6442_65;
  wire  T_6442_66;
  wire  T_6442_67;
  wire  T_6442_68;
  wire  T_6442_69;
  wire  T_6442_70;
  wire  T_6442_71;
  wire  T_6442_72;
  wire  T_6442_73;
  wire  T_6442_74;
  wire  T_6442_75;
  wire  T_6442_76;
  wire  T_6442_77;
  wire  T_6442_78;
  wire  T_6442_79;
  wire  T_6442_80;
  wire  T_6442_81;
  wire  T_6442_82;
  wire  T_6442_83;
  wire  T_6442_84;
  wire  T_6442_85;
  wire  T_6442_86;
  wire  T_6442_87;
  wire  T_6442_88;
  wire  T_6442_89;
  wire  T_6442_90;
  wire  T_6442_91;
  wire  T_6442_92;
  wire  T_6442_93;
  wire  T_6442_94;
  wire  T_6442_95;
  wire  T_6442_96;
  wire  T_6442_97;
  wire  T_6442_98;
  wire  T_6442_99;
  wire  T_6442_100;
  wire  T_6442_101;
  wire  T_6442_102;
  wire  T_6442_103;
  wire  T_6442_104;
  wire  T_6442_105;
  wire  T_6442_106;
  wire  T_6442_107;
  wire  T_6442_108;
  wire  T_6442_109;
  wire  T_6442_110;
  wire  T_6442_111;
  wire  T_6442_112;
  wire  T_6442_113;
  wire  T_6442_114;
  wire  T_6442_115;
  wire  T_6442_116;
  wire  T_6442_117;
  wire  T_6442_118;
  wire  T_6442_119;
  wire  T_6442_120;
  wire  T_6442_121;
  wire  T_6442_122;
  wire  T_6442_123;
  wire  T_6442_124;
  wire  T_6442_125;
  wire  T_6442_126;
  wire  T_6442_127;
  wire  T_6576;
  wire  T_6583;
  wire  T_6587;
  wire  T_6591;
  wire  T_6598;
  wire  T_6602;
  wire  T_6606;
  wire  T_6631;
  wire  T_6638;
  wire  T_6642;
  wire  T_6646;
  wire  T_6653;
  wire  T_6657;
  wire  T_6661;
  wire  T_6686;
  wire  T_6690;
  wire  T_6694;
  wire  T_6698;
  wire  T_6702;
  wire  T_6706;
  wire  T_6710;
  wire  T_6714;
  wire  T_6718;
  wire  T_6722;
  wire  T_6726;
  wire  T_6730;
  wire  T_6734;
  wire  T_6738;
  wire  T_6742;
  wire  T_6746;
  wire  T_6798;
  wire  T_6802;
  wire  T_6806;
  wire  T_6810;
  wire  T_6814;
  wire  T_6818;
  wire  T_6822;
  wire  T_6826;
  wire  T_6830;
  wire  T_6834;
  wire  T_6838;
  wire  T_6842;
  wire  T_6846;
  wire  T_6850;
  wire  T_6854;
  wire  T_6858;
  wire  T_6862;
  wire  T_6866;
  wire  T_6870;
  wire  T_6874;
  wire  T_7138_0;
  wire  T_7138_1;
  wire  T_7138_2;
  wire  T_7138_3;
  wire  T_7138_4;
  wire  T_7138_5;
  wire  T_7138_6;
  wire  T_7138_7;
  wire  T_7138_8;
  wire  T_7138_9;
  wire  T_7138_10;
  wire  T_7138_11;
  wire  T_7138_12;
  wire  T_7138_13;
  wire  T_7138_14;
  wire  T_7138_15;
  wire  T_7138_16;
  wire  T_7138_17;
  wire  T_7138_18;
  wire  T_7138_19;
  wire  T_7138_20;
  wire  T_7138_21;
  wire  T_7138_22;
  wire  T_7138_23;
  wire  T_7138_24;
  wire  T_7138_25;
  wire  T_7138_26;
  wire  T_7138_27;
  wire  T_7138_28;
  wire  T_7138_29;
  wire  T_7138_30;
  wire  T_7138_31;
  wire  T_7138_32;
  wire  T_7138_33;
  wire  T_7138_34;
  wire  T_7138_35;
  wire  T_7138_36;
  wire  T_7138_37;
  wire  T_7138_38;
  wire  T_7138_39;
  wire  T_7138_40;
  wire  T_7138_41;
  wire  T_7138_42;
  wire  T_7138_43;
  wire  T_7138_44;
  wire  T_7138_45;
  wire  T_7138_46;
  wire  T_7138_47;
  wire  T_7138_48;
  wire  T_7138_49;
  wire  T_7138_50;
  wire  T_7138_51;
  wire  T_7138_52;
  wire  T_7138_53;
  wire  T_7138_54;
  wire  T_7138_55;
  wire  T_7138_56;
  wire  T_7138_57;
  wire  T_7138_58;
  wire  T_7138_59;
  wire  T_7138_60;
  wire  T_7138_61;
  wire  T_7138_62;
  wire  T_7138_63;
  wire  T_7138_64;
  wire  T_7138_65;
  wire  T_7138_66;
  wire  T_7138_67;
  wire  T_7138_68;
  wire  T_7138_69;
  wire  T_7138_70;
  wire  T_7138_71;
  wire  T_7138_72;
  wire  T_7138_73;
  wire  T_7138_74;
  wire  T_7138_75;
  wire  T_7138_76;
  wire  T_7138_77;
  wire  T_7138_78;
  wire  T_7138_79;
  wire  T_7138_80;
  wire  T_7138_81;
  wire  T_7138_82;
  wire  T_7138_83;
  wire  T_7138_84;
  wire  T_7138_85;
  wire  T_7138_86;
  wire  T_7138_87;
  wire  T_7138_88;
  wire  T_7138_89;
  wire  T_7138_90;
  wire  T_7138_91;
  wire  T_7138_92;
  wire  T_7138_93;
  wire  T_7138_94;
  wire  T_7138_95;
  wire  T_7138_96;
  wire  T_7138_97;
  wire  T_7138_98;
  wire  T_7138_99;
  wire  T_7138_100;
  wire  T_7138_101;
  wire  T_7138_102;
  wire  T_7138_103;
  wire  T_7138_104;
  wire  T_7138_105;
  wire  T_7138_106;
  wire  T_7138_107;
  wire  T_7138_108;
  wire  T_7138_109;
  wire  T_7138_110;
  wire  T_7138_111;
  wire  T_7138_112;
  wire  T_7138_113;
  wire  T_7138_114;
  wire  T_7138_115;
  wire  T_7138_116;
  wire  T_7138_117;
  wire  T_7138_118;
  wire  T_7138_119;
  wire  T_7138_120;
  wire  T_7138_121;
  wire  T_7138_122;
  wire  T_7138_123;
  wire  T_7138_124;
  wire  T_7138_125;
  wire  T_7138_126;
  wire  T_7138_127;
  wire  T_7269;
  wire  T_7270;
  wire  T_7271;
  wire  T_7272;
  wire  T_7273;
  wire  T_7274;
  wire  T_7275;
  wire [1:0] T_7279;
  wire [2:0] T_7280;
  wire [1:0] T_7281;
  wire [1:0] T_7282;
  wire [3:0] T_7283;
  wire [6:0] T_7284;
  wire  T_7285;
  wire  T_7286;
  wire  T_7287;
  wire  T_7288;
  wire  T_7289;
  wire  T_7290;
  wire  T_7291;
  wire [1:0] T_7295;
  wire [2:0] T_7296;
  wire [1:0] T_7297;
  wire [1:0] T_7298;
  wire [3:0] T_7299;
  wire [6:0] T_7300;
  wire  GEN_0;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_58;
  wire  GEN_59;
  wire  GEN_60;
  wire  GEN_61;
  wire  GEN_62;
  wire  GEN_63;
  wire  GEN_64;
  wire  GEN_65;
  wire  GEN_66;
  wire  GEN_67;
  wire  GEN_68;
  wire  GEN_69;
  wire  GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  wire  GEN_73;
  wire  GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  GEN_77;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_85;
  wire  GEN_86;
  wire  GEN_87;
  wire  GEN_88;
  wire  GEN_89;
  wire  GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_95;
  wire  GEN_96;
  wire  GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire  GEN_106;
  wire  GEN_107;
  wire  GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire  GEN_113;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  GEN_117;
  wire  GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire  GEN_128;
  wire  GEN_129;
  wire  GEN_130;
  wire  GEN_131;
  wire  GEN_132;
  wire  GEN_133;
  wire  GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire  GEN_140;
  wire  GEN_141;
  wire  GEN_142;
  wire  GEN_143;
  wire  GEN_144;
  wire  GEN_145;
  wire  GEN_146;
  wire  GEN_147;
  wire  GEN_148;
  wire  GEN_1;
  wire  GEN_149;
  wire  GEN_150;
  wire  GEN_151;
  wire  GEN_152;
  wire  GEN_153;
  wire  GEN_154;
  wire  GEN_155;
  wire  GEN_156;
  wire  GEN_157;
  wire  GEN_158;
  wire  GEN_159;
  wire  GEN_160;
  wire  GEN_161;
  wire  GEN_162;
  wire  GEN_163;
  wire  GEN_164;
  wire  GEN_165;
  wire  GEN_166;
  wire  GEN_167;
  wire  GEN_168;
  wire  GEN_169;
  wire  GEN_170;
  wire  GEN_171;
  wire  GEN_172;
  wire  GEN_173;
  wire  GEN_174;
  wire  GEN_175;
  wire  GEN_176;
  wire  GEN_177;
  wire  GEN_178;
  wire  GEN_179;
  wire  GEN_180;
  wire  GEN_181;
  wire  GEN_182;
  wire  GEN_183;
  wire  GEN_184;
  wire  GEN_185;
  wire  GEN_186;
  wire  GEN_187;
  wire  GEN_188;
  wire  GEN_189;
  wire  GEN_190;
  wire  GEN_191;
  wire  GEN_192;
  wire  GEN_193;
  wire  GEN_194;
  wire  GEN_195;
  wire  GEN_196;
  wire  GEN_197;
  wire  GEN_198;
  wire  GEN_199;
  wire  GEN_200;
  wire  GEN_201;
  wire  GEN_202;
  wire  GEN_203;
  wire  GEN_204;
  wire  GEN_205;
  wire  GEN_206;
  wire  GEN_207;
  wire  GEN_208;
  wire  GEN_209;
  wire  GEN_210;
  wire  GEN_211;
  wire  GEN_212;
  wire  GEN_213;
  wire  GEN_214;
  wire  GEN_215;
  wire  GEN_216;
  wire  GEN_217;
  wire  GEN_218;
  wire  GEN_219;
  wire  GEN_220;
  wire  GEN_221;
  wire  GEN_222;
  wire  GEN_223;
  wire  GEN_224;
  wire  GEN_225;
  wire  GEN_226;
  wire  GEN_227;
  wire  GEN_228;
  wire  GEN_229;
  wire  GEN_230;
  wire  GEN_231;
  wire  GEN_232;
  wire  GEN_233;
  wire  GEN_234;
  wire  GEN_235;
  wire  GEN_236;
  wire  GEN_237;
  wire  GEN_238;
  wire  GEN_239;
  wire  GEN_240;
  wire  GEN_241;
  wire  GEN_242;
  wire  GEN_243;
  wire  GEN_244;
  wire  GEN_245;
  wire  GEN_246;
  wire  GEN_247;
  wire  GEN_248;
  wire  GEN_249;
  wire  GEN_250;
  wire  GEN_251;
  wire  GEN_252;
  wire  GEN_253;
  wire  GEN_254;
  wire  GEN_255;
  wire  GEN_256;
  wire  GEN_257;
  wire  GEN_258;
  wire  GEN_259;
  wire  GEN_260;
  wire  GEN_261;
  wire  GEN_262;
  wire  GEN_263;
  wire  GEN_264;
  wire  GEN_265;
  wire  GEN_266;
  wire  GEN_267;
  wire  GEN_268;
  wire  GEN_269;
  wire  GEN_270;
  wire  GEN_271;
  wire  GEN_272;
  wire  GEN_273;
  wire  GEN_274;
  wire  GEN_275;
  wire  T_7303;
  wire  GEN_2;
  wire  GEN_276;
  wire  GEN_277;
  wire  GEN_278;
  wire  GEN_279;
  wire  GEN_280;
  wire  GEN_281;
  wire  GEN_282;
  wire  GEN_283;
  wire  GEN_284;
  wire  GEN_285;
  wire  GEN_286;
  wire  GEN_287;
  wire  GEN_288;
  wire  GEN_289;
  wire  GEN_290;
  wire  GEN_291;
  wire  GEN_292;
  wire  GEN_293;
  wire  GEN_294;
  wire  GEN_295;
  wire  GEN_296;
  wire  GEN_297;
  wire  GEN_298;
  wire  GEN_299;
  wire  GEN_300;
  wire  GEN_301;
  wire  GEN_302;
  wire  GEN_303;
  wire  GEN_304;
  wire  GEN_305;
  wire  GEN_306;
  wire  GEN_307;
  wire  GEN_308;
  wire  GEN_309;
  wire  GEN_310;
  wire  GEN_311;
  wire  GEN_312;
  wire  GEN_313;
  wire  GEN_314;
  wire  GEN_315;
  wire  GEN_316;
  wire  GEN_317;
  wire  GEN_318;
  wire  GEN_319;
  wire  GEN_320;
  wire  GEN_321;
  wire  GEN_322;
  wire  GEN_323;
  wire  GEN_324;
  wire  GEN_325;
  wire  GEN_326;
  wire  GEN_327;
  wire  GEN_328;
  wire  GEN_329;
  wire  GEN_330;
  wire  GEN_331;
  wire  GEN_332;
  wire  GEN_333;
  wire  GEN_334;
  wire  GEN_335;
  wire  GEN_336;
  wire  GEN_337;
  wire  GEN_338;
  wire  GEN_339;
  wire  GEN_340;
  wire  GEN_341;
  wire  GEN_342;
  wire  GEN_343;
  wire  GEN_344;
  wire  GEN_345;
  wire  GEN_346;
  wire  GEN_347;
  wire  GEN_348;
  wire  GEN_349;
  wire  GEN_350;
  wire  GEN_351;
  wire  GEN_352;
  wire  GEN_353;
  wire  GEN_354;
  wire  GEN_355;
  wire  GEN_356;
  wire  GEN_357;
  wire  GEN_358;
  wire  GEN_359;
  wire  GEN_360;
  wire  GEN_361;
  wire  GEN_362;
  wire  GEN_363;
  wire  GEN_364;
  wire  GEN_365;
  wire  GEN_366;
  wire  GEN_367;
  wire  GEN_368;
  wire  GEN_369;
  wire  GEN_370;
  wire  GEN_371;
  wire  GEN_372;
  wire  GEN_373;
  wire  GEN_374;
  wire  GEN_375;
  wire  GEN_376;
  wire  GEN_377;
  wire  GEN_378;
  wire  GEN_379;
  wire  GEN_380;
  wire  GEN_381;
  wire  GEN_382;
  wire  GEN_383;
  wire  GEN_384;
  wire  GEN_385;
  wire  GEN_386;
  wire  GEN_387;
  wire  GEN_388;
  wire  GEN_389;
  wire  GEN_390;
  wire  GEN_391;
  wire  GEN_392;
  wire  GEN_393;
  wire  GEN_394;
  wire  GEN_395;
  wire  GEN_396;
  wire  GEN_397;
  wire  GEN_398;
  wire  GEN_399;
  wire  GEN_400;
  wire  GEN_401;
  wire  GEN_402;
  wire  GEN_3;
  wire  GEN_403;
  wire  GEN_404;
  wire  GEN_405;
  wire  GEN_406;
  wire  GEN_407;
  wire  GEN_408;
  wire  GEN_409;
  wire  GEN_410;
  wire  GEN_411;
  wire  GEN_412;
  wire  GEN_413;
  wire  GEN_414;
  wire  GEN_415;
  wire  GEN_416;
  wire  GEN_417;
  wire  GEN_418;
  wire  GEN_419;
  wire  GEN_420;
  wire  GEN_421;
  wire  GEN_422;
  wire  GEN_423;
  wire  GEN_424;
  wire  GEN_425;
  wire  GEN_426;
  wire  GEN_427;
  wire  GEN_428;
  wire  GEN_429;
  wire  GEN_430;
  wire  GEN_431;
  wire  GEN_432;
  wire  GEN_433;
  wire  GEN_434;
  wire  GEN_435;
  wire  GEN_436;
  wire  GEN_437;
  wire  GEN_438;
  wire  GEN_439;
  wire  GEN_440;
  wire  GEN_441;
  wire  GEN_442;
  wire  GEN_443;
  wire  GEN_444;
  wire  GEN_445;
  wire  GEN_446;
  wire  GEN_447;
  wire  GEN_448;
  wire  GEN_449;
  wire  GEN_450;
  wire  GEN_451;
  wire  GEN_452;
  wire  GEN_453;
  wire  GEN_454;
  wire  GEN_455;
  wire  GEN_456;
  wire  GEN_457;
  wire  GEN_458;
  wire  GEN_459;
  wire  GEN_460;
  wire  GEN_461;
  wire  GEN_462;
  wire  GEN_463;
  wire  GEN_464;
  wire  GEN_465;
  wire  GEN_466;
  wire  GEN_467;
  wire  GEN_468;
  wire  GEN_469;
  wire  GEN_470;
  wire  GEN_471;
  wire  GEN_472;
  wire  GEN_473;
  wire  GEN_474;
  wire  GEN_475;
  wire  GEN_476;
  wire  GEN_477;
  wire  GEN_478;
  wire  GEN_479;
  wire  GEN_480;
  wire  GEN_481;
  wire  GEN_482;
  wire  GEN_483;
  wire  GEN_484;
  wire  GEN_485;
  wire  GEN_486;
  wire  GEN_487;
  wire  GEN_488;
  wire  GEN_489;
  wire  GEN_490;
  wire  GEN_491;
  wire  GEN_492;
  wire  GEN_493;
  wire  GEN_494;
  wire  GEN_495;
  wire  GEN_496;
  wire  GEN_497;
  wire  GEN_498;
  wire  GEN_499;
  wire  GEN_500;
  wire  GEN_501;
  wire  GEN_502;
  wire  GEN_503;
  wire  GEN_504;
  wire  GEN_505;
  wire  GEN_506;
  wire  GEN_507;
  wire  GEN_508;
  wire  GEN_509;
  wire  GEN_510;
  wire  GEN_511;
  wire  GEN_512;
  wire  GEN_513;
  wire  GEN_514;
  wire  GEN_515;
  wire  GEN_516;
  wire  GEN_517;
  wire  GEN_518;
  wire  GEN_519;
  wire  GEN_520;
  wire  GEN_521;
  wire  GEN_522;
  wire  GEN_523;
  wire  GEN_524;
  wire  GEN_525;
  wire  GEN_526;
  wire  GEN_527;
  wire  GEN_528;
  wire  GEN_529;
  wire  T_7306;
  wire  T_7307;
  wire  T_7308;
  wire  T_7309;
  wire  T_7310;
  wire [127:0] T_7312;
  wire [1:0] T_7313;
  wire [1:0] T_7314;
  wire [3:0] T_7315;
  wire [1:0] T_7316;
  wire [1:0] T_7317;
  wire [3:0] T_7318;
  wire [7:0] T_7319;
  wire [1:0] T_7320;
  wire [3:0] T_7322;
  wire [7:0] T_7326;
  wire [15:0] T_7327;
  wire [1:0] T_7328;
  wire [1:0] T_7329;
  wire [3:0] T_7330;
  wire [1:0] T_7331;
  wire [1:0] T_7332;
  wire [3:0] T_7333;
  wire [7:0] T_7334;
  wire [1:0] T_7335;
  wire [3:0] T_7337;
  wire [7:0] T_7341;
  wire [15:0] T_7342;
  wire [31:0] T_7343;
  wire [1:0] T_7344;
  wire [1:0] T_7345;
  wire [3:0] T_7346;
  wire [1:0] T_7347;
  wire [1:0] T_7348;
  wire [3:0] T_7349;
  wire [7:0] T_7350;
  wire [1:0] T_7351;
  wire [1:0] T_7352;
  wire [3:0] T_7353;
  wire [1:0] T_7354;
  wire [1:0] T_7355;
  wire [3:0] T_7356;
  wire [7:0] T_7357;
  wire [15:0] T_7358;
  wire [31:0] T_7374;
  wire [63:0] T_7375;
  wire [1:0] T_7376;
  wire [1:0] T_7377;
  wire [3:0] T_7378;
  wire [1:0] T_7379;
  wire [1:0] T_7380;
  wire [3:0] T_7381;
  wire [7:0] T_7382;
  wire [1:0] T_7383;
  wire [1:0] T_7384;
  wire [3:0] T_7385;
  wire [1:0] T_7386;
  wire [1:0] T_7387;
  wire [3:0] T_7388;
  wire [7:0] T_7389;
  wire [15:0] T_7390;
  wire [1:0] T_7391;
  wire [1:0] T_7392;
  wire [3:0] T_7393;
  wire [7:0] T_7397;
  wire [15:0] T_7405;
  wire [31:0] T_7406;
  wire [63:0] T_7438;
  wire [127:0] T_7439;
  wire [127:0] T_7440;
  wire [127:0] T_7442;
  wire [1:0] T_7443;
  wire [1:0] T_7444;
  wire [3:0] T_7445;
  wire [1:0] T_7446;
  wire [1:0] T_7447;
  wire [3:0] T_7448;
  wire [7:0] T_7449;
  wire [1:0] T_7450;
  wire [3:0] T_7452;
  wire [7:0] T_7456;
  wire [15:0] T_7457;
  wire [1:0] T_7458;
  wire [1:0] T_7459;
  wire [3:0] T_7460;
  wire [1:0] T_7461;
  wire [1:0] T_7462;
  wire [3:0] T_7463;
  wire [7:0] T_7464;
  wire [1:0] T_7465;
  wire [3:0] T_7467;
  wire [7:0] T_7471;
  wire [15:0] T_7472;
  wire [31:0] T_7473;
  wire [1:0] T_7474;
  wire [1:0] T_7475;
  wire [3:0] T_7476;
  wire [1:0] T_7477;
  wire [1:0] T_7478;
  wire [3:0] T_7479;
  wire [7:0] T_7480;
  wire [1:0] T_7481;
  wire [1:0] T_7482;
  wire [3:0] T_7483;
  wire [1:0] T_7484;
  wire [1:0] T_7485;
  wire [3:0] T_7486;
  wire [7:0] T_7487;
  wire [15:0] T_7488;
  wire [31:0] T_7504;
  wire [63:0] T_7505;
  wire [1:0] T_7506;
  wire [1:0] T_7507;
  wire [3:0] T_7508;
  wire [1:0] T_7509;
  wire [1:0] T_7510;
  wire [3:0] T_7511;
  wire [7:0] T_7512;
  wire [1:0] T_7513;
  wire [1:0] T_7514;
  wire [3:0] T_7515;
  wire [1:0] T_7516;
  wire [1:0] T_7517;
  wire [3:0] T_7518;
  wire [7:0] T_7519;
  wire [15:0] T_7520;
  wire [1:0] T_7521;
  wire [1:0] T_7522;
  wire [3:0] T_7523;
  wire [7:0] T_7527;
  wire [15:0] T_7535;
  wire [31:0] T_7536;
  wire [63:0] T_7568;
  wire [127:0] T_7569;
  wire [127:0] T_7570;
  wire  T_7571;
  wire  T_7572;
  wire  T_7573;
  wire  T_7574;
  wire  T_7577;
  wire  T_7578;
  wire  T_7580;
  wire  T_7581;
  wire  T_7582;
  wire  T_7583;
  wire  T_7584;
  wire  T_7587;
  wire  T_7588;
  wire  T_7590;
  wire  T_7613;
  wire  T_7614;
  wire  T_7620;
  wire  T_7623;
  wire  T_7624;
  wire  T_7630;
  wire  T_7633;
  wire  T_7634;
  wire  T_7640;
  wire  T_7643;
  wire  T_7644;
  wire  T_7650;
  wire  T_7653;
  wire  T_7654;
  wire  T_7660;
  wire  T_7663;
  wire  T_7664;
  wire  T_7670;
  wire  T_7693;
  wire  T_7694;
  wire  T_7700;
  wire  T_7703;
  wire  T_7704;
  wire  T_7710;
  wire  T_7713;
  wire  T_7714;
  wire  T_7720;
  wire  T_7723;
  wire  T_7724;
  wire  T_7730;
  wire  T_7733;
  wire  T_7734;
  wire  T_7740;
  wire  T_7743;
  wire  T_7744;
  wire  T_7750;
  wire  T_7893;
  wire  T_7894;
  wire  T_7900;
  wire  T_7903;
  wire  T_7904;
  wire  T_7910;
  wire  T_7933;
  wire  T_7934;
  wire  T_7940;
  wire  T_7943;
  wire  T_7944;
  wire  T_7950;
  wire  T_7953;
  wire  T_7954;
  wire  T_7960;
  wire  T_7963;
  wire  T_7964;
  wire  T_7970;
  wire  T_7973;
  wire  T_7974;
  wire  T_7980;
  wire  T_7983;
  wire  T_7984;
  wire  T_7990;
  wire  T_8013;
  wire  T_8014;
  wire  T_8020;
  wire  T_8023;
  wire  T_8024;
  wire  T_8030;
  wire  T_8033;
  wire  T_8034;
  wire  T_8040;
  wire  T_8043;
  wire  T_8044;
  wire  T_8050;
  wire  T_8053;
  wire  T_8054;
  wire  T_8060;
  wire  T_8063;
  wire  T_8064;
  wire  T_8070;
  wire  T_8213;
  wire  T_8214;
  wire  T_8220;
  wire  T_8223;
  wire  T_8224;
  wire  T_8230;
  wire  T_8233;
  wire  T_8234;
  wire  T_8240;
  wire  T_8243;
  wire  T_8244;
  wire  T_8250;
  wire  T_8253;
  wire  T_8254;
  wire  T_8260;
  wire  T_8263;
  wire  T_8264;
  wire  T_8270;
  wire  T_8273;
  wire  T_8274;
  wire  T_8280;
  wire  T_8283;
  wire  T_8284;
  wire  T_8290;
  wire  T_8293;
  wire  T_8294;
  wire  T_8300;
  wire  T_8303;
  wire  T_8304;
  wire  T_8310;
  wire  T_8313;
  wire  T_8314;
  wire  T_8320;
  wire  T_8323;
  wire  T_8324;
  wire  T_8330;
  wire  T_8333;
  wire  T_8334;
  wire  T_8340;
  wire  T_8343;
  wire  T_8344;
  wire  T_8350;
  wire  T_8353;
  wire  T_8354;
  wire  T_8360;
  wire  T_8363;
  wire  T_8364;
  wire  T_8370;
  wire  T_8373;
  wire  T_8374;
  wire  T_8380;
  wire  T_8383;
  wire  T_8384;
  wire  T_8390;
  wire  T_8393;
  wire  T_8394;
  wire  T_8400;
  wire  T_8403;
  wire  T_8404;
  wire  T_8410;
  wire  T_8413;
  wire  T_8414;
  wire  T_8420;
  wire  T_8423;
  wire  T_8424;
  wire  T_8430;
  wire  T_8433;
  wire  T_8434;
  wire  T_8440;
  wire  T_8443;
  wire  T_8444;
  wire  T_8450;
  wire  T_8453;
  wire  T_8454;
  wire  T_8460;
  wire  T_8463;
  wire  T_8464;
  wire  T_8470;
  wire  T_8473;
  wire  T_8474;
  wire  T_8480;
  wire  T_8483;
  wire  T_8484;
  wire  T_8490;
  wire  T_8493;
  wire  T_8494;
  wire  T_8500;
  wire  T_8503;
  wire  T_8504;
  wire  T_8510;
  wire  T_8513;
  wire  T_8514;
  wire  T_8520;
  wire  T_8523;
  wire  T_8524;
  wire  T_8530;
  wire  T_8853;
  wire  T_8854;
  wire  T_8860;
  wire  T_8863;
  wire  T_8864;
  wire  T_8870;
  wire  T_8873;
  wire  T_8874;
  wire  T_8880;
  wire  T_8883;
  wire  T_8884;
  wire  T_8890;
  wire  T_8893;
  wire  T_8894;
  wire  T_8900;
  wire  T_8903;
  wire  T_8904;
  wire  T_8910;
  wire  T_8913;
  wire  T_8914;
  wire  T_8920;
  wire  T_8923;
  wire  T_8924;
  wire  T_8930;
  wire  T_8933;
  wire  T_8934;
  wire  T_8940;
  wire  T_8943;
  wire  T_8944;
  wire  T_8950;
  wire  T_8953;
  wire  T_8954;
  wire  T_8960;
  wire  T_8963;
  wire  T_8964;
  wire  T_8970;
  wire  T_8973;
  wire  T_8974;
  wire  T_8980;
  wire  T_8983;
  wire  T_8984;
  wire  T_8990;
  wire  T_8993;
  wire  T_8994;
  wire  T_9000;
  wire  T_9003;
  wire  T_9004;
  wire  T_9010;
  wire  T_9013;
  wire  T_9014;
  wire  T_9020;
  wire  T_9023;
  wire  T_9024;
  wire  T_9030;
  wire  T_9033;
  wire  T_9034;
  wire  T_9040;
  wire  T_9043;
  wire  T_9044;
  wire  T_9050;
  wire  T_9053;
  wire  T_9054;
  wire  T_9060;
  wire  T_9063;
  wire  T_9064;
  wire  T_9070;
  wire  T_9073;
  wire  T_9074;
  wire  T_9080;
  wire  T_9083;
  wire  T_9084;
  wire  T_9090;
  wire  T_9093;
  wire  T_9094;
  wire  T_9100;
  wire  T_9103;
  wire  T_9104;
  wire  T_9110;
  wire  T_9113;
  wire  T_9114;
  wire  T_9120;
  wire  T_9123;
  wire  T_9124;
  wire  T_9130;
  wire  T_9133;
  wire  T_9134;
  wire  T_9140;
  wire  T_9143;
  wire  T_9144;
  wire  T_9150;
  wire  T_9153;
  wire  T_9154;
  wire  T_9160;
  wire  T_9163;
  wire  T_9164;
  wire  T_9170;
  wire  T_9173;
  wire  T_9174;
  wire  T_9180;
  wire  T_9183;
  wire  T_9184;
  wire  T_9190;
  wire  T_9193;
  wire  T_9194;
  wire  T_9200;
  wire  T_9203;
  wire  T_9204;
  wire  T_9210;
  wire  T_9213;
  wire  T_9214;
  wire  T_9220;
  wire  T_9223;
  wire  T_9224;
  wire  T_9230;
  wire  T_9233;
  wire  T_9234;
  wire  T_9240;
  wire  T_9243;
  wire  T_9244;
  wire  T_9250;
  wire  T_10462_0;
  wire  T_10462_1;
  wire  T_10462_2;
  wire  T_10462_3;
  wire  T_10462_4;
  wire  T_10462_5;
  wire  T_10462_6;
  wire  T_10462_7;
  wire  T_10462_8;
  wire  T_10462_9;
  wire  T_10462_10;
  wire  T_10462_11;
  wire  T_10462_12;
  wire  T_10462_13;
  wire  T_10462_14;
  wire  T_10462_15;
  wire  T_10462_16;
  wire  T_10462_17;
  wire  T_10462_18;
  wire  T_10462_19;
  wire  T_10462_20;
  wire  T_10462_21;
  wire  T_10462_22;
  wire  T_10462_23;
  wire  T_10462_24;
  wire  T_10462_25;
  wire  T_10462_26;
  wire  T_10462_27;
  wire  T_10462_28;
  wire  T_10462_29;
  wire  T_10462_30;
  wire  T_10462_31;
  wire  T_10462_32;
  wire  T_10462_33;
  wire  T_10462_34;
  wire  T_10462_35;
  wire  T_10462_36;
  wire  T_10462_37;
  wire  T_10462_38;
  wire  T_10462_39;
  wire  T_10462_40;
  wire  T_10462_41;
  wire  T_10462_42;
  wire  T_10462_43;
  wire  T_10462_44;
  wire  T_10462_45;
  wire  T_10462_46;
  wire  T_10462_47;
  wire  T_10462_48;
  wire  T_10462_49;
  wire  T_10462_50;
  wire  T_10462_51;
  wire  T_10462_52;
  wire  T_10462_53;
  wire  T_10462_54;
  wire  T_10462_55;
  wire  T_10462_56;
  wire  T_10462_57;
  wire  T_10462_58;
  wire  T_10462_59;
  wire  T_10462_60;
  wire  T_10462_61;
  wire  T_10462_62;
  wire  T_10462_63;
  wire  T_10462_64;
  wire  T_10462_65;
  wire  T_10462_66;
  wire  T_10462_67;
  wire  T_10462_68;
  wire  T_10462_69;
  wire  T_10462_70;
  wire  T_10462_71;
  wire  T_10462_72;
  wire  T_10462_73;
  wire  T_10462_74;
  wire  T_10462_75;
  wire  T_10462_76;
  wire  T_10462_77;
  wire  T_10462_78;
  wire  T_10462_79;
  wire  T_10462_80;
  wire  T_10462_81;
  wire  T_10462_82;
  wire  T_10462_83;
  wire  T_10462_84;
  wire  T_10462_85;
  wire  T_10462_86;
  wire  T_10462_87;
  wire  T_10462_88;
  wire  T_10462_89;
  wire  T_10462_90;
  wire  T_10462_91;
  wire  T_10462_92;
  wire  T_10462_93;
  wire  T_10462_94;
  wire  T_10462_95;
  wire  T_10462_96;
  wire  T_10462_97;
  wire  T_10462_98;
  wire  T_10462_99;
  wire  T_10462_100;
  wire  T_10462_101;
  wire  T_10462_102;
  wire  T_10462_103;
  wire  T_10462_104;
  wire  T_10462_105;
  wire  T_10462_106;
  wire  T_10462_107;
  wire  T_10462_108;
  wire  T_10462_109;
  wire  T_10462_110;
  wire  T_10462_111;
  wire  T_10462_112;
  wire  T_10462_113;
  wire  T_10462_114;
  wire  T_10462_115;
  wire  T_10462_116;
  wire  T_10462_117;
  wire  T_10462_118;
  wire  T_10462_119;
  wire  T_10462_120;
  wire  T_10462_121;
  wire  T_10462_122;
  wire  T_10462_123;
  wire  T_10462_124;
  wire  T_10462_125;
  wire  T_10462_126;
  wire  T_10462_127;
  wire [31:0] T_10725_0;
  wire [31:0] T_10725_1;
  wire [31:0] T_10725_2;
  wire [31:0] T_10725_3;
  wire [31:0] T_10725_4;
  wire [31:0] T_10725_5;
  wire [31:0] T_10725_6;
  wire [31:0] T_10725_7;
  wire [31:0] T_10725_8;
  wire [31:0] T_10725_9;
  wire [31:0] T_10725_10;
  wire [31:0] T_10725_11;
  wire [31:0] T_10725_12;
  wire [31:0] T_10725_13;
  wire [31:0] T_10725_14;
  wire [31:0] T_10725_15;
  wire [31:0] T_10725_16;
  wire [31:0] T_10725_17;
  wire [31:0] T_10725_18;
  wire [31:0] T_10725_19;
  wire [31:0] T_10725_20;
  wire [31:0] T_10725_21;
  wire [31:0] T_10725_22;
  wire [31:0] T_10725_23;
  wire [31:0] T_10725_24;
  wire [31:0] T_10725_25;
  wire [31:0] T_10725_26;
  wire [31:0] T_10725_27;
  wire [31:0] T_10725_28;
  wire [31:0] T_10725_29;
  wire [31:0] T_10725_30;
  wire [31:0] T_10725_31;
  wire [31:0] T_10725_32;
  wire [31:0] T_10725_33;
  wire [31:0] T_10725_34;
  wire [31:0] T_10725_35;
  wire [31:0] T_10725_36;
  wire [31:0] T_10725_37;
  wire [31:0] T_10725_38;
  wire [31:0] T_10725_39;
  wire [31:0] T_10725_40;
  wire [31:0] T_10725_41;
  wire [31:0] T_10725_42;
  wire [31:0] T_10725_43;
  wire [31:0] T_10725_44;
  wire [31:0] T_10725_45;
  wire [31:0] T_10725_46;
  wire [31:0] T_10725_47;
  wire [31:0] T_10725_48;
  wire [31:0] T_10725_49;
  wire [31:0] T_10725_50;
  wire [31:0] T_10725_51;
  wire [31:0] T_10725_52;
  wire [31:0] T_10725_53;
  wire [31:0] T_10725_54;
  wire [31:0] T_10725_55;
  wire [31:0] T_10725_56;
  wire [31:0] T_10725_57;
  wire [31:0] T_10725_58;
  wire [31:0] T_10725_59;
  wire [31:0] T_10725_60;
  wire [31:0] T_10725_61;
  wire [31:0] T_10725_62;
  wire [31:0] T_10725_63;
  wire [31:0] T_10725_64;
  wire [31:0] T_10725_65;
  wire [31:0] T_10725_66;
  wire [31:0] T_10725_67;
  wire [31:0] T_10725_68;
  wire [31:0] T_10725_69;
  wire [31:0] T_10725_70;
  wire [31:0] T_10725_71;
  wire [31:0] T_10725_72;
  wire [31:0] T_10725_73;
  wire [31:0] T_10725_74;
  wire [31:0] T_10725_75;
  wire [31:0] T_10725_76;
  wire [31:0] T_10725_77;
  wire [31:0] T_10725_78;
  wire [31:0] T_10725_79;
  wire [31:0] T_10725_80;
  wire [31:0] T_10725_81;
  wire [31:0] T_10725_82;
  wire [31:0] T_10725_83;
  wire [31:0] T_10725_84;
  wire [31:0] T_10725_85;
  wire [31:0] T_10725_86;
  wire [31:0] T_10725_87;
  wire [31:0] T_10725_88;
  wire [31:0] T_10725_89;
  wire [31:0] T_10725_90;
  wire [31:0] T_10725_91;
  wire [31:0] T_10725_92;
  wire [31:0] T_10725_93;
  wire [31:0] T_10725_94;
  wire [31:0] T_10725_95;
  wire [31:0] T_10725_96;
  wire [31:0] T_10725_97;
  wire [31:0] T_10725_98;
  wire [31:0] T_10725_99;
  wire [31:0] T_10725_100;
  wire [31:0] T_10725_101;
  wire [31:0] T_10725_102;
  wire [31:0] T_10725_103;
  wire [31:0] T_10725_104;
  wire [31:0] T_10725_105;
  wire [31:0] T_10725_106;
  wire [31:0] T_10725_107;
  wire [31:0] T_10725_108;
  wire [31:0] T_10725_109;
  wire [31:0] T_10725_110;
  wire [31:0] T_10725_111;
  wire [31:0] T_10725_112;
  wire [31:0] T_10725_113;
  wire [31:0] T_10725_114;
  wire [31:0] T_10725_115;
  wire [31:0] T_10725_116;
  wire [31:0] T_10725_117;
  wire [31:0] T_10725_118;
  wire [31:0] T_10725_119;
  wire [31:0] T_10725_120;
  wire [31:0] T_10725_121;
  wire [31:0] T_10725_122;
  wire [31:0] T_10725_123;
  wire [31:0] T_10725_124;
  wire [31:0] T_10725_125;
  wire [31:0] T_10725_126;
  wire [31:0] T_10725_127;
  wire  GEN_4;
  wire  GEN_530;
  wire  GEN_531;
  wire  GEN_532;
  wire  GEN_533;
  wire  GEN_534;
  wire  GEN_535;
  wire  GEN_536;
  wire  GEN_537;
  wire  GEN_538;
  wire  GEN_539;
  wire  GEN_540;
  wire  GEN_541;
  wire  GEN_542;
  wire  GEN_543;
  wire  GEN_544;
  wire  GEN_545;
  wire  GEN_546;
  wire  GEN_547;
  wire  GEN_548;
  wire  GEN_549;
  wire  GEN_550;
  wire  GEN_551;
  wire  GEN_552;
  wire  GEN_553;
  wire  GEN_554;
  wire  GEN_555;
  wire  GEN_556;
  wire  GEN_557;
  wire  GEN_558;
  wire  GEN_559;
  wire  GEN_560;
  wire  GEN_561;
  wire  GEN_562;
  wire  GEN_563;
  wire  GEN_564;
  wire  GEN_565;
  wire  GEN_566;
  wire  GEN_567;
  wire  GEN_568;
  wire  GEN_569;
  wire  GEN_570;
  wire  GEN_571;
  wire  GEN_572;
  wire  GEN_573;
  wire  GEN_574;
  wire  GEN_575;
  wire  GEN_576;
  wire  GEN_577;
  wire  GEN_578;
  wire  GEN_579;
  wire  GEN_580;
  wire  GEN_581;
  wire  GEN_582;
  wire  GEN_583;
  wire  GEN_584;
  wire  GEN_585;
  wire  GEN_586;
  wire  GEN_587;
  wire  GEN_588;
  wire  GEN_589;
  wire  GEN_590;
  wire  GEN_591;
  wire  GEN_592;
  wire  GEN_593;
  wire  GEN_594;
  wire  GEN_595;
  wire  GEN_596;
  wire  GEN_597;
  wire  GEN_598;
  wire  GEN_599;
  wire  GEN_600;
  wire  GEN_601;
  wire  GEN_602;
  wire  GEN_603;
  wire  GEN_604;
  wire  GEN_605;
  wire  GEN_606;
  wire  GEN_607;
  wire  GEN_608;
  wire  GEN_609;
  wire  GEN_610;
  wire  GEN_611;
  wire  GEN_612;
  wire  GEN_613;
  wire  GEN_614;
  wire  GEN_615;
  wire  GEN_616;
  wire  GEN_617;
  wire  GEN_618;
  wire  GEN_619;
  wire  GEN_620;
  wire  GEN_621;
  wire  GEN_622;
  wire  GEN_623;
  wire  GEN_624;
  wire  GEN_625;
  wire  GEN_626;
  wire  GEN_627;
  wire  GEN_628;
  wire  GEN_629;
  wire  GEN_630;
  wire  GEN_631;
  wire  GEN_632;
  wire  GEN_633;
  wire  GEN_634;
  wire  GEN_635;
  wire  GEN_636;
  wire  GEN_637;
  wire  GEN_638;
  wire  GEN_639;
  wire  GEN_640;
  wire  GEN_641;
  wire  GEN_642;
  wire  GEN_643;
  wire  GEN_644;
  wire  GEN_645;
  wire  GEN_646;
  wire  GEN_647;
  wire  GEN_648;
  wire  GEN_649;
  wire  GEN_650;
  wire  GEN_651;
  wire  GEN_652;
  wire  GEN_653;
  wire  GEN_654;
  wire  GEN_655;
  wire  GEN_656;
  wire [31:0] GEN_5;
  wire [31:0] GEN_657;
  wire [31:0] GEN_658;
  wire [31:0] GEN_659;
  wire [31:0] GEN_660;
  wire [31:0] GEN_661;
  wire [31:0] GEN_662;
  wire [31:0] GEN_663;
  wire [31:0] GEN_664;
  wire [31:0] GEN_665;
  wire [31:0] GEN_666;
  wire [31:0] GEN_667;
  wire [31:0] GEN_668;
  wire [31:0] GEN_669;
  wire [31:0] GEN_670;
  wire [31:0] GEN_671;
  wire [31:0] GEN_672;
  wire [31:0] GEN_673;
  wire [31:0] GEN_674;
  wire [31:0] GEN_675;
  wire [31:0] GEN_676;
  wire [31:0] GEN_677;
  wire [31:0] GEN_678;
  wire [31:0] GEN_679;
  wire [31:0] GEN_680;
  wire [31:0] GEN_681;
  wire [31:0] GEN_682;
  wire [31:0] GEN_683;
  wire [31:0] GEN_684;
  wire [31:0] GEN_685;
  wire [31:0] GEN_686;
  wire [31:0] GEN_687;
  wire [31:0] GEN_688;
  wire [31:0] GEN_689;
  wire [31:0] GEN_690;
  wire [31:0] GEN_691;
  wire [31:0] GEN_692;
  wire [31:0] GEN_693;
  wire [31:0] GEN_694;
  wire [31:0] GEN_695;
  wire [31:0] GEN_696;
  wire [31:0] GEN_697;
  wire [31:0] GEN_698;
  wire [31:0] GEN_699;
  wire [31:0] GEN_700;
  wire [31:0] GEN_701;
  wire [31:0] GEN_702;
  wire [31:0] GEN_703;
  wire [31:0] GEN_704;
  wire [31:0] GEN_705;
  wire [31:0] GEN_706;
  wire [31:0] GEN_707;
  wire [31:0] GEN_708;
  wire [31:0] GEN_709;
  wire [31:0] GEN_710;
  wire [31:0] GEN_711;
  wire [31:0] GEN_712;
  wire [31:0] GEN_713;
  wire [31:0] GEN_714;
  wire [31:0] GEN_715;
  wire [31:0] GEN_716;
  wire [31:0] GEN_717;
  wire [31:0] GEN_718;
  wire [31:0] GEN_719;
  wire [31:0] GEN_720;
  wire [31:0] GEN_721;
  wire [31:0] GEN_722;
  wire [31:0] GEN_723;
  wire [31:0] GEN_724;
  wire [31:0] GEN_725;
  wire [31:0] GEN_726;
  wire [31:0] GEN_727;
  wire [31:0] GEN_728;
  wire [31:0] GEN_729;
  wire [31:0] GEN_730;
  wire [31:0] GEN_731;
  wire [31:0] GEN_732;
  wire [31:0] GEN_733;
  wire [31:0] GEN_734;
  wire [31:0] GEN_735;
  wire [31:0] GEN_736;
  wire [31:0] GEN_737;
  wire [31:0] GEN_738;
  wire [31:0] GEN_739;
  wire [31:0] GEN_740;
  wire [31:0] GEN_741;
  wire [31:0] GEN_742;
  wire [31:0] GEN_743;
  wire [31:0] GEN_744;
  wire [31:0] GEN_745;
  wire [31:0] GEN_746;
  wire [31:0] GEN_747;
  wire [31:0] GEN_748;
  wire [31:0] GEN_749;
  wire [31:0] GEN_750;
  wire [31:0] GEN_751;
  wire [31:0] GEN_752;
  wire [31:0] GEN_753;
  wire [31:0] GEN_754;
  wire [31:0] GEN_755;
  wire [31:0] GEN_756;
  wire [31:0] GEN_757;
  wire [31:0] GEN_758;
  wire [31:0] GEN_759;
  wire [31:0] GEN_760;
  wire [31:0] GEN_761;
  wire [31:0] GEN_762;
  wire [31:0] GEN_763;
  wire [31:0] GEN_764;
  wire [31:0] GEN_765;
  wire [31:0] GEN_766;
  wire [31:0] GEN_767;
  wire [31:0] GEN_768;
  wire [31:0] GEN_769;
  wire [31:0] GEN_770;
  wire [31:0] GEN_771;
  wire [31:0] GEN_772;
  wire [31:0] GEN_773;
  wire [31:0] GEN_774;
  wire [31:0] GEN_775;
  wire [31:0] GEN_776;
  wire [31:0] GEN_777;
  wire [31:0] GEN_778;
  wire [31:0] GEN_779;
  wire [31:0] GEN_780;
  wire [31:0] GEN_781;
  wire [31:0] GEN_782;
  wire [31:0] GEN_783;
  wire [31:0] T_10858;
  wire [1:0] T_10859;
  wire [4:0] T_10861;
  wire [2:0] T_10862;
  wire [2:0] T_10873_opcode;
  wire [1:0] T_10873_param;
  wire [2:0] T_10873_size;
  wire [4:0] T_10873_source;
  wire  T_10873_sink;
  wire [1:0] T_10873_addr_lo;
  wire [31:0] T_10873_data;
  wire  T_10873_error;
  wire [2:0] GEN_784 = 3'b0;
  reg [31:0] GEN_808;
  wire [1:0] GEN_785 = 2'b0;
  reg [31:0] GEN_809;
  wire [2:0] GEN_786 = 3'b0;
  reg [31:0] GEN_810;
  wire [4:0] GEN_787 = 5'b0;
  reg [31:0] GEN_811;
  wire [28:0] GEN_788 = 29'b0;
  reg [31:0] GEN_812;
  wire [3:0] GEN_789 = 4'b0;
  reg [31:0] GEN_813;
  wire [31:0] GEN_790 = 32'b0;
  reg [31:0] GEN_814;
  wire  GEN_791 = 1'b0;
  reg [31:0] GEN_815;
  sirv_rtc rtc (
    .clock(rtc_clock),
    .reset(rtc_reset),
    .io_regs_cfg_write_valid(rtc_io_regs_cfg_write_valid),
    .io_regs_cfg_write_bits(rtc_io_regs_cfg_write_bits),
    .io_regs_cfg_read(rtc_io_regs_cfg_read),
    .io_regs_countLo_write_valid(rtc_io_regs_countLo_write_valid),
    .io_regs_countLo_write_bits(rtc_io_regs_countLo_write_bits),
    .io_regs_countLo_read(rtc_io_regs_countLo_read),
    .io_regs_countHi_write_valid(rtc_io_regs_countHi_write_valid),
    .io_regs_countHi_write_bits(rtc_io_regs_countHi_write_bits),
    .io_regs_countHi_read(rtc_io_regs_countHi_read),
    .io_regs_s_write_valid(rtc_io_regs_s_write_valid),
    .io_regs_s_write_bits(rtc_io_regs_s_write_bits),
    .io_regs_s_read(rtc_io_regs_s_read),
    .io_regs_cmp_0_write_valid(rtc_io_regs_cmp_0_write_valid),
    .io_regs_cmp_0_write_bits(rtc_io_regs_cmp_0_write_bits),
    .io_regs_cmp_0_read(rtc_io_regs_cmp_0_read),
    .io_regs_feed_write_valid(rtc_io_regs_feed_write_valid),
    .io_regs_feed_write_bits(rtc_io_regs_feed_write_bits),
    .io_regs_feed_read(rtc_io_regs_feed_read),
    .io_regs_key_write_valid(rtc_io_regs_key_write_valid),
    .io_regs_key_write_bits(rtc_io_regs_key_write_bits),
    .io_regs_key_read(rtc_io_regs_key_read),
    .io_ip_0(rtc_io_ip_0)
  );
  sirv_pmu u_sirv_pmu (
    .clock(pmu_clock),
    .reset(pmu_reset),
    .io_wakeup_awakeup(pmu_io_wakeup_awakeup),
    .io_wakeup_dwakeup(pmu_io_wakeup_dwakeup),
    .io_wakeup_rtc(pmu_io_wakeup_rtc),
    .io_wakeup_reset(pmu_io_wakeup_reset),
    .io_control_hfclkrst(pmu_io_control_hfclkrst),
    .io_control_corerst(pmu_io_control_corerst),
    .io_control_reserved1(pmu_io_control_reserved1),
    .io_control_vddpaden(pmu_io_control_vddpaden),
    .io_control_reserved0(pmu_io_control_reserved0),
    .io_regs_ie_write_valid(pmu_io_regs_ie_write_valid),
    .io_regs_ie_write_bits(pmu_io_regs_ie_write_bits),
    .io_regs_ie_read(pmu_io_regs_ie_read),
    .io_regs_cause_write_valid(pmu_io_regs_cause_write_valid),
    .io_regs_cause_write_bits(pmu_io_regs_cause_write_bits),
    .io_regs_cause_read(pmu_io_regs_cause_read),
    .io_regs_sleep_write_valid(pmu_io_regs_sleep_write_valid),
    .io_regs_sleep_write_bits(pmu_io_regs_sleep_write_bits),
    .io_regs_sleep_read(pmu_io_regs_sleep_read),
    .io_regs_key_write_valid(pmu_io_regs_key_write_valid),
    .io_regs_key_write_bits(pmu_io_regs_key_write_bits),
    .io_regs_key_read(pmu_io_regs_key_read),
    .io_regs_wakeupProgram_0_write_valid(pmu_io_regs_wakeupProgram_0_write_valid),
    .io_regs_wakeupProgram_0_write_bits(pmu_io_regs_wakeupProgram_0_write_bits),
    .io_regs_wakeupProgram_0_read(pmu_io_regs_wakeupProgram_0_read),
    .io_regs_wakeupProgram_1_write_valid(pmu_io_regs_wakeupProgram_1_write_valid),
    .io_regs_wakeupProgram_1_write_bits(pmu_io_regs_wakeupProgram_1_write_bits),
    .io_regs_wakeupProgram_1_read(pmu_io_regs_wakeupProgram_1_read),
    .io_regs_wakeupProgram_2_write_valid(pmu_io_regs_wakeupProgram_2_write_valid),
    .io_regs_wakeupProgram_2_write_bits(pmu_io_regs_wakeupProgram_2_write_bits),
    .io_regs_wakeupProgram_2_read(pmu_io_regs_wakeupProgram_2_read),
    .io_regs_wakeupProgram_3_write_valid(pmu_io_regs_wakeupProgram_3_write_valid),
    .io_regs_wakeupProgram_3_write_bits(pmu_io_regs_wakeupProgram_3_write_bits),
    .io_regs_wakeupProgram_3_read(pmu_io_regs_wakeupProgram_3_read),
    .io_regs_wakeupProgram_4_write_valid(pmu_io_regs_wakeupProgram_4_write_valid),
    .io_regs_wakeupProgram_4_write_bits(pmu_io_regs_wakeupProgram_4_write_bits),
    .io_regs_wakeupProgram_4_read(pmu_io_regs_wakeupProgram_4_read),
    .io_regs_wakeupProgram_5_write_valid(pmu_io_regs_wakeupProgram_5_write_valid),
    .io_regs_wakeupProgram_5_write_bits(pmu_io_regs_wakeupProgram_5_write_bits),
    .io_regs_wakeupProgram_5_read(pmu_io_regs_wakeupProgram_5_read),
    .io_regs_wakeupProgram_6_write_valid(pmu_io_regs_wakeupProgram_6_write_valid),
    .io_regs_wakeupProgram_6_write_bits(pmu_io_regs_wakeupProgram_6_write_bits),
    .io_regs_wakeupProgram_6_read(pmu_io_regs_wakeupProgram_6_read),
    .io_regs_wakeupProgram_7_write_valid(pmu_io_regs_wakeupProgram_7_write_valid),
    .io_regs_wakeupProgram_7_write_bits(pmu_io_regs_wakeupProgram_7_write_bits),
    .io_regs_wakeupProgram_7_read(pmu_io_regs_wakeupProgram_7_read),
    .io_regs_sleepProgram_0_write_valid(pmu_io_regs_sleepProgram_0_write_valid),
    .io_regs_sleepProgram_0_write_bits(pmu_io_regs_sleepProgram_0_write_bits),
    .io_regs_sleepProgram_0_read(pmu_io_regs_sleepProgram_0_read),
    .io_regs_sleepProgram_1_write_valid(pmu_io_regs_sleepProgram_1_write_valid),
    .io_regs_sleepProgram_1_write_bits(pmu_io_regs_sleepProgram_1_write_bits),
    .io_regs_sleepProgram_1_read(pmu_io_regs_sleepProgram_1_read),
    .io_regs_sleepProgram_2_write_valid(pmu_io_regs_sleepProgram_2_write_valid),
    .io_regs_sleepProgram_2_write_bits(pmu_io_regs_sleepProgram_2_write_bits),
    .io_regs_sleepProgram_2_read(pmu_io_regs_sleepProgram_2_read),
    .io_regs_sleepProgram_3_write_valid(pmu_io_regs_sleepProgram_3_write_valid),
    .io_regs_sleepProgram_3_write_bits(pmu_io_regs_sleepProgram_3_write_bits),
    .io_regs_sleepProgram_3_read(pmu_io_regs_sleepProgram_3_read),
    .io_regs_sleepProgram_4_write_valid(pmu_io_regs_sleepProgram_4_write_valid),
    .io_regs_sleepProgram_4_write_bits(pmu_io_regs_sleepProgram_4_write_bits),
    .io_regs_sleepProgram_4_read(pmu_io_regs_sleepProgram_4_read),
    .io_regs_sleepProgram_5_write_valid(pmu_io_regs_sleepProgram_5_write_valid),
    .io_regs_sleepProgram_5_write_bits(pmu_io_regs_sleepProgram_5_write_bits),
    .io_regs_sleepProgram_5_read(pmu_io_regs_sleepProgram_5_read),
    .io_regs_sleepProgram_6_write_valid(pmu_io_regs_sleepProgram_6_write_valid),
    .io_regs_sleepProgram_6_write_bits(pmu_io_regs_sleepProgram_6_write_bits),
    .io_regs_sleepProgram_6_read(pmu_io_regs_sleepProgram_6_read),
    .io_regs_sleepProgram_7_write_valid(pmu_io_regs_sleepProgram_7_write_valid),
    .io_regs_sleepProgram_7_write_bits(pmu_io_regs_sleepProgram_7_write_bits),
    .io_regs_sleepProgram_7_read(pmu_io_regs_sleepProgram_7_read),
    .io_resetCauses_wdogrst(pmu_io_resetCauses_wdogrst),
    .io_resetCauses_erst(pmu_io_resetCauses_erst),
    .io_resetCauses_porrst(pmu_io_resetCauses_porrst)
  );
  sirv_wdog wdog (
    .clock(wdog_clock),
    .reset(wdog_reset),
    .io_regs_cfg_write_valid(wdog_io_regs_cfg_write_valid),
    .io_regs_cfg_write_bits(wdog_io_regs_cfg_write_bits),
    .io_regs_cfg_read(wdog_io_regs_cfg_read),
    .io_regs_countLo_write_valid(wdog_io_regs_countLo_write_valid),
    .io_regs_countLo_write_bits(wdog_io_regs_countLo_write_bits),
    .io_regs_countLo_read(wdog_io_regs_countLo_read),
    .io_regs_countHi_write_valid(wdog_io_regs_countHi_write_valid),
    .io_regs_countHi_write_bits(wdog_io_regs_countHi_write_bits),
    .io_regs_countHi_read(wdog_io_regs_countHi_read),
    .io_regs_s_write_valid(wdog_io_regs_s_write_valid),
    .io_regs_s_write_bits(wdog_io_regs_s_write_bits),
    .io_regs_s_read(wdog_io_regs_s_read),
    .io_regs_cmp_0_write_valid(wdog_io_regs_cmp_0_write_valid),
    .io_regs_cmp_0_write_bits(wdog_io_regs_cmp_0_write_bits),
    .io_regs_cmp_0_read(wdog_io_regs_cmp_0_read),
    .io_regs_feed_write_valid(wdog_io_regs_feed_write_valid),
    .io_regs_feed_write_bits(wdog_io_regs_feed_write_bits),
    .io_regs_feed_read(wdog_io_regs_feed_read),
    .io_regs_key_write_valid(wdog_io_regs_key_write_valid),
    .io_regs_key_write_bits(wdog_io_regs_key_write_bits),
    .io_regs_key_read(wdog_io_regs_key_read),
    .io_ip_0(wdog_io_ip_0),
    .io_corerst(wdog_io_corerst),
    .io_rst(wdog_io_rst)
  );
  sirv_queue u_queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_read(Queue_1_io_enq_bits_read),
    .io_enq_bits_index(Queue_1_io_enq_bits_index),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_mask(Queue_1_io_enq_bits_mask),
    .io_enq_bits_extra(Queue_1_io_enq_bits_extra),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_read(Queue_1_io_deq_bits_read),
    .io_deq_bits_index(Queue_1_io_deq_bits_index),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_mask(Queue_1_io_deq_bits_mask),
    .io_deq_bits_extra(Queue_1_io_deq_bits_extra),
    .io_count(Queue_1_io_count)
  );
  assign io_interrupts_0_0 = wdog_io_ip_0;
  assign io_interrupts_0_1 = rtc_io_ip_0;
  assign io_in_0_a_ready = T_953_ready;
  assign io_in_0_b_valid = 1'h0;
  assign io_in_0_b_bits_opcode = GEN_784;
  assign io_in_0_b_bits_param = GEN_785;
  assign io_in_0_b_bits_size = GEN_786;
  assign io_in_0_b_bits_source = GEN_787;
  assign io_in_0_b_bits_address = GEN_788;
  assign io_in_0_b_bits_mask = GEN_789;
  assign io_in_0_b_bits_data = GEN_790;
  assign io_in_0_c_ready = 1'h1;
  assign io_in_0_d_valid = T_992_valid;
  assign io_in_0_d_bits_opcode = {{2'd0}, T_992_bits_read};
  assign io_in_0_d_bits_param = T_10873_param;
  assign io_in_0_d_bits_size = T_10873_size;
  assign io_in_0_d_bits_source = T_10873_source;
  assign io_in_0_d_bits_sink = T_10873_sink;
  assign io_in_0_d_bits_addr_lo = T_10873_addr_lo;
  assign io_in_0_d_bits_data = T_992_bits_data;
  assign io_in_0_d_bits_error = T_10873_error;
  assign io_in_0_e_ready = 1'h1;
  // assign io_lfclk = io_lfextclk;
   CLKBUFUHDV4 u_buf_io_lfclk( 
    .Z(io_lfclk     ),
    .I(io_lfextclk  )
 );

  // In DFT mode the internal generated reset siganls should be disabled
  assign io_moff_hfclkrst = test_mode ? erst : pmu_io_control_hfclkrst;
  assign io_moff_corerst  = test_mode ? erst : pmu_io_control_corerst;
  assign io_wdog_rst      = test_mode ? erst : wdog_io_rst;

        //Bob: This reserved1 signal is actually the padrst signal used in hifive board
  assign io_pmu_padrst = test_mode ? 1'b1 : pmu_io_control_reserved1;

  // In DFT mode the power control siganls should be disabled
  assign io_pmu_vddpaden  = test_mode ? 1'b1 : pmu_io_control_vddpaden;

  assign rtc_clock = clock;
  assign rtc_reset = reset;
  assign rtc_io_regs_cfg_write_valid = T_3904;
  assign rtc_io_regs_cfg_write_bits = T_2505;
  assign rtc_io_regs_countLo_write_valid = T_3824;
  assign rtc_io_regs_countLo_write_bits = T_2505;
  assign rtc_io_regs_countHi_write_valid = T_4264;
  assign rtc_io_regs_countHi_write_bits = T_2505;
  assign rtc_io_regs_s_write_valid = T_2704;
  assign rtc_io_regs_s_write_bits = T_2505;
  assign rtc_io_regs_cmp_0_write_valid = T_2624;
  assign rtc_io_regs_cmp_0_write_bits = T_2505;
  assign rtc_io_regs_feed_write_valid = T_3384;
  assign rtc_io_regs_feed_write_bits = T_2505;
  assign rtc_io_regs_key_write_valid = T_4064;
  assign rtc_io_regs_key_write_bits = T_2505;
  assign pmu_clock = clock;
  assign pmu_reset = reset;
  assign pmu_io_wakeup_awakeup = 1'h0;
  assign pmu_io_wakeup_dwakeup = io_pmu_dwakeup;
  assign pmu_io_wakeup_rtc = rtc_io_ip_0;
  assign pmu_io_wakeup_reset = GEN_791;
  assign pmu_io_regs_ie_write_valid = T_3744;
  assign pmu_io_regs_ie_write_bits = T_3745;
  assign pmu_io_regs_cause_write_valid = T_3504;
  assign pmu_io_regs_cause_write_bits = T_2505;
  assign pmu_io_regs_sleep_write_valid = T_4184;
  assign pmu_io_regs_sleep_write_bits = T_2505;
  assign pmu_io_regs_key_write_valid = T_4464;
  assign pmu_io_regs_key_write_bits = T_2505;
  assign pmu_io_regs_wakeupProgram_0_write_valid = T_3344;
  assign pmu_io_regs_wakeupProgram_0_write_bits = T_2505;
  assign pmu_io_regs_wakeupProgram_1_write_valid = T_3024;
  assign pmu_io_regs_wakeupProgram_1_write_bits = T_2505;
  assign pmu_io_regs_wakeupProgram_2_write_valid = T_3664;
  assign pmu_io_regs_wakeupProgram_2_write_bits = T_2505;
  assign pmu_io_regs_wakeupProgram_3_write_valid = T_3864;
  assign pmu_io_regs_wakeupProgram_3_write_bits = T_2505;
  assign pmu_io_regs_wakeupProgram_4_write_valid = T_4424;
  assign pmu_io_regs_wakeupProgram_4_write_bits = T_2505;
  assign pmu_io_regs_wakeupProgram_5_write_valid = T_2504;
  assign pmu_io_regs_wakeupProgram_5_write_bits = T_2505;
  assign pmu_io_regs_wakeupProgram_6_write_valid = T_2944;
  assign pmu_io_regs_wakeupProgram_6_write_bits = T_2505;
  assign pmu_io_regs_wakeupProgram_7_write_valid = T_3464;
  assign pmu_io_regs_wakeupProgram_7_write_bits = T_2505;
  assign pmu_io_regs_sleepProgram_0_write_valid = T_3944;
  assign pmu_io_regs_sleepProgram_0_write_bits = T_2505;
  assign pmu_io_regs_sleepProgram_1_write_valid = T_3144;
  assign pmu_io_regs_sleepProgram_1_write_bits = T_2505;
  assign pmu_io_regs_sleepProgram_2_write_valid = T_2824;
  assign pmu_io_regs_sleepProgram_2_write_bits = T_2505;
  assign pmu_io_regs_sleepProgram_3_write_valid = T_4144;
  assign pmu_io_regs_sleepProgram_3_write_bits = T_2505;
  assign pmu_io_regs_sleepProgram_4_write_valid = T_3544;
  assign pmu_io_regs_sleepProgram_4_write_bits = T_2505;
  assign pmu_io_regs_sleepProgram_5_write_valid = T_3064;
  assign pmu_io_regs_sleepProgram_5_write_bits = T_2505;
  assign pmu_io_regs_sleepProgram_6_write_valid = T_2784;
  assign pmu_io_regs_sleepProgram_6_write_bits = T_2505;
  assign pmu_io_regs_sleepProgram_7_write_valid = T_4344;
  assign pmu_io_regs_sleepProgram_7_write_bits = T_2505;
  assign pmu_io_resetCauses_wdogrst = io_resetCauses_wdogrst;
  assign pmu_io_resetCauses_erst = io_resetCauses_erst;
  assign pmu_io_resetCauses_porrst = io_resetCauses_porrst;
  assign wdog_clock = clock;
  assign wdog_reset = reset;
  assign wdog_io_regs_cfg_write_valid = T_2544;
  assign wdog_io_regs_cfg_write_bits = T_2505;
  assign wdog_io_regs_countLo_write_valid = T_3184;
  assign wdog_io_regs_countLo_write_bits = T_2505;
  assign wdog_io_regs_countHi_write_valid = T_3704;
  assign wdog_io_regs_countHi_write_bits = T_2505;
  assign wdog_io_regs_s_write_valid = T_4304;
  assign wdog_io_regs_s_write_bits = T_4105;
  assign wdog_io_regs_cmp_0_write_valid = T_4104;
  assign wdog_io_regs_cmp_0_write_bits = T_4105;
  assign wdog_io_regs_feed_write_valid = T_2864;
  assign wdog_io_regs_feed_write_bits = T_2505;
  assign wdog_io_regs_key_write_valid = T_3584;
  assign wdog_io_regs_key_write_bits = T_2505;
  assign wdog_io_corerst = pmu_io_control_corerst;
  assign T_953_ready = T_7307;
  assign T_953_valid = io_in_0_a_valid;
  assign T_953_bits_read = T_970;
  assign T_953_bits_index = T_971[9:0];
  assign T_953_bits_data = io_in_0_a_bits_data;
  assign T_953_bits_mask = io_in_0_a_bits_mask;
  assign T_953_bits_extra = T_974;
  assign T_970 = io_in_0_a_bits_opcode == 3'h4;
  assign T_971 = io_in_0_a_bits_address[28:2];
  assign T_972 = io_in_0_a_bits_address[1:0];
  assign T_973 = {T_972,io_in_0_a_bits_source};
  assign T_974 = {T_973,io_in_0_a_bits_size};
  assign T_992_ready = io_in_0_d_ready;
  assign T_992_valid = T_7310;
  assign T_992_bits_read = Queue_1_io_deq_bits_read;
  assign T_992_bits_data = T_10858;
  assign T_992_bits_extra = Queue_1_io_deq_bits_extra;
  assign T_1028_ready = Queue_1_io_enq_ready;
  assign T_1028_valid = T_7308;
  assign T_1028_bits_read = T_953_bits_read;
  assign T_1028_bits_index = T_953_bits_index;
  assign T_1028_bits_data = T_953_bits_data;
  assign T_1028_bits_mask = T_953_bits_mask;
  assign T_1028_bits_extra = T_953_bits_extra;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = T_1028_valid;
  assign Queue_1_io_enq_bits_read = T_1028_bits_read;
  assign Queue_1_io_enq_bits_index = T_1028_bits_index;
  assign Queue_1_io_enq_bits_data = T_1028_bits_data;
  assign Queue_1_io_enq_bits_mask = T_1028_bits_mask;
  assign Queue_1_io_enq_bits_extra = T_1028_bits_extra;
  assign Queue_1_io_deq_ready = T_7309;
  assign T_1310 = T_1028_bits_index ^ 10'h45;
  assign T_1311 = T_1310 & 10'h380;
  assign T_1313 = T_1311 == 10'h0;
  assign T_1314 = Queue_1_io_deq_bits_index ^ 10'h45;
  assign T_1315 = T_1314 & 10'h380;
  assign T_1317 = T_1315 == 10'h0;
  assign T_1320 = T_1028_bits_index & 10'h380;
  assign T_1322 = T_1320 == 10'h0;
  assign T_1323 = Queue_1_io_deq_bits_index;
  assign T_1324 = T_1323 & 10'h380;
  assign T_1326 = T_1324 == 10'h0;
  assign T_1328 = T_1028_bits_index ^ 10'h2a;
  assign T_1329 = T_1328 & 10'h380;
  assign T_1331 = T_1329 == 10'h0;
  assign T_1332 = Queue_1_io_deq_bits_index ^ 10'h2a;
  assign T_1333 = T_1332 & 10'h380;
  assign T_1335 = T_1333 == 10'h0;
  assign T_1337 = T_1028_bits_index ^ 10'h18;
  assign T_1338 = T_1337 & 10'h380;
  assign T_1340 = T_1338 == 10'h0;
  assign T_1341 = Queue_1_io_deq_bits_index ^ 10'h18;
  assign T_1342 = T_1341 & 10'h380;
  assign T_1344 = T_1342 == 10'h0;
  assign T_1346 = T_1028_bits_index ^ 10'h25;
  assign T_1347 = T_1346 & 10'h380;
  assign T_1349 = T_1347 == 10'h0;
  assign T_1350 = Queue_1_io_deq_bits_index ^ 10'h25;
  assign T_1351 = T_1350 & 10'h380;
  assign T_1353 = T_1351 == 10'h0;
  assign T_1355 = T_1028_bits_index ^ 10'h14;
  assign T_1356 = T_1355 & 10'h380;
  assign T_1358 = T_1356 == 10'h0;
  assign T_1359 = Queue_1_io_deq_bits_index ^ 10'h14;
  assign T_1360 = T_1359 & 10'h380;
  assign T_1362 = T_1360 == 10'h0;
  assign T_1364 = T_1028_bits_index ^ 10'h2e;
  assign T_1365 = T_1364 & 10'h380;
  assign T_1367 = T_1365 == 10'h0;
  assign T_1368 = Queue_1_io_deq_bits_index ^ 10'h2e;
  assign T_1369 = T_1368 & 10'h380;
  assign T_1371 = T_1369 == 10'h0;
  assign T_1373 = T_1028_bits_index ^ 10'h4e;
  assign T_1374 = T_1373 & 10'h380;
  assign T_1376 = T_1374 == 10'h0;
  assign T_1377 = Queue_1_io_deq_bits_index ^ 10'h4e;
  assign T_1378 = T_1377 & 10'h380;
  assign T_1380 = T_1378 == 10'h0;
  assign T_1382 = T_1028_bits_index ^ 10'h4a;
  assign T_1383 = T_1382 & 10'h380;
  assign T_1385 = T_1383 == 10'h0;
  assign T_1386 = Queue_1_io_deq_bits_index ^ 10'h4a;
  assign T_1387 = T_1386 & 10'h380;
  assign T_1389 = T_1387 == 10'h0;
  assign T_1391 = T_1028_bits_index ^ 10'h6;
  assign T_1392 = T_1391 & 10'h380;
  assign T_1394 = T_1392 == 10'h0;
  assign T_1395 = Queue_1_io_deq_bits_index ^ 10'h6;
  assign T_1396 = T_1395 & 10'h380;
  assign T_1398 = T_1396 == 10'h0;
  assign T_1400 = T_1028_bits_index ^ 10'h26;
  assign T_1401 = T_1400 & 10'h380;
  assign T_1403 = T_1401 == 10'h0;
  assign T_1404 = Queue_1_io_deq_bits_index ^ 10'h26;
  assign T_1405 = T_1404 & 10'h380;
  assign T_1407 = T_1405 == 10'h0;
  assign T_1409 = T_1028_bits_index ^ 10'h46;
  assign T_1410 = T_1409 & 10'h380;
  assign T_1412 = T_1410 == 10'h0;
  assign T_1413 = Queue_1_io_deq_bits_index ^ 10'h46;
  assign T_1414 = T_1413 & 10'h380;
  assign T_1416 = T_1414 == 10'h0;
  assign T_1418 = T_1028_bits_index ^ 10'h21;
  assign T_1419 = T_1418 & 10'h380;
  assign T_1421 = T_1419 == 10'h0;
  assign T_1422 = Queue_1_io_deq_bits_index ^ 10'h21;
  assign T_1423 = T_1422 & 10'h380;
  assign T_1425 = T_1423 == 10'h0;
  assign T_1427 = T_1028_bits_index ^ 10'h41;
  assign T_1428 = T_1427 & 10'h380;
  assign T_1430 = T_1428 == 10'h0;
  assign T_1431 = Queue_1_io_deq_bits_index ^ 10'h41;
  assign T_1432 = T_1431 & 10'h380;
  assign T_1434 = T_1432 == 10'h0;
  assign T_1436 = T_1028_bits_index ^ 10'h4d;
  assign T_1437 = T_1436 & 10'h380;
  assign T_1439 = T_1437 == 10'h0;
  assign T_1440 = Queue_1_io_deq_bits_index ^ 10'h4d;
  assign T_1441 = T_1440 & 10'h380;
  assign T_1443 = T_1441 == 10'h0;
  assign T_1445 = T_1028_bits_index ^ 10'h29;
  assign T_1446 = T_1445 & 10'h380;
  assign T_1448 = T_1446 == 10'h0;
  assign T_1449 = Queue_1_io_deq_bits_index ^ 10'h29;
  assign T_1450 = T_1449 & 10'h380;
  assign T_1452 = T_1450 == 10'h0;
  assign T_1454 = T_1028_bits_index ^ 10'h49;
  assign T_1455 = T_1454 & 10'h380;
  assign T_1457 = T_1455 == 10'h0;
  assign T_1458 = Queue_1_io_deq_bits_index ^ 10'h49;
  assign T_1459 = T_1458 & 10'h380;
  assign T_1461 = T_1459 == 10'h0;
  assign T_1463 = T_1028_bits_index ^ 10'h2;
  assign T_1464 = T_1463 & 10'h380;
  assign T_1466 = T_1464 == 10'h0;
  assign T_1467 = Queue_1_io_deq_bits_index ^ 10'h2;
  assign T_1468 = T_1467 & 10'h380;
  assign T_1470 = T_1468 == 10'h0;
  assign T_1472 = T_1028_bits_index ^ 10'h20;
  assign T_1473 = T_1472 & 10'h380;
  assign T_1475 = T_1473 == 10'h0;
  assign T_1476 = Queue_1_io_deq_bits_index ^ 10'h20;
  assign T_1477 = T_1476 & 10'h380;
  assign T_1479 = T_1477 == 10'h0;
  assign T_1481 = T_1028_bits_index ^ 10'h22;
  assign T_1482 = T_1481 & 10'h380;
  assign T_1484 = T_1482 == 10'h0;
  assign T_1485 = Queue_1_io_deq_bits_index ^ 10'h22;
  assign T_1486 = T_1485 & 10'h380;
  assign T_1488 = T_1486 == 10'h0;
  assign T_1490 = T_1028_bits_index ^ 10'h2d;
  assign T_1491 = T_1490 & 10'h380;
  assign T_1493 = T_1491 == 10'h0;
  assign T_1494 = Queue_1_io_deq_bits_index ^ 10'h2d;
  assign T_1495 = T_1494 & 10'h380;
  assign T_1497 = T_1495 == 10'h0;
  assign T_1499 = T_1028_bits_index ^ 10'h40;
  assign T_1500 = T_1499 & 10'h380;
  assign T_1502 = T_1500 == 10'h0;
  assign T_1503 = Queue_1_io_deq_bits_index ^ 10'h40;
  assign T_1504 = T_1503 & 10'h380;
  assign T_1506 = T_1504 == 10'h0;
  assign T_1508 = T_1028_bits_index ^ 10'h16;
  assign T_1509 = T_1508 & 10'h380;
  assign T_1511 = T_1509 == 10'h0;
  assign T_1512 = Queue_1_io_deq_bits_index ^ 10'h16;
  assign T_1513 = T_1512 & 10'h380;
  assign T_1515 = T_1513 == 10'h0;
  assign T_1517 = T_1028_bits_index ^ 10'h2c;
  assign T_1518 = T_1517 & 10'h380;
  assign T_1520 = T_1518 == 10'h0;
  assign T_1521 = Queue_1_io_deq_bits_index ^ 10'h2c;
  assign T_1522 = T_1521 & 10'h380;
  assign T_1524 = T_1522 == 10'h0;
  assign T_1526 = T_1028_bits_index ^ 10'h47;
  assign T_1527 = T_1526 & 10'h380;
  assign T_1529 = T_1527 == 10'h0;
  assign T_1530 = Queue_1_io_deq_bits_index ^ 10'h47;
  assign T_1531 = T_1530 & 10'h380;
  assign T_1533 = T_1531 == 10'h0;
  assign T_1535 = T_1028_bits_index ^ 10'h51;
  assign T_1536 = T_1535 & 10'h380;
  assign T_1538 = T_1536 == 10'h0;
  assign T_1539 = Queue_1_io_deq_bits_index ^ 10'h51;
  assign T_1540 = T_1539 & 10'h380;
  assign T_1542 = T_1540 == 10'h0;
  assign T_1544 = T_1028_bits_index ^ 10'h4c;
  assign T_1545 = T_1544 & 10'h380;
  assign T_1547 = T_1545 == 10'h0;
  assign T_1548 = Queue_1_io_deq_bits_index ^ 10'h4c;
  assign T_1549 = T_1548 & 10'h380;
  assign T_1551 = T_1549 == 10'h0;
  assign T_1553 = T_1028_bits_index ^ 10'h7;
  assign T_1554 = T_1553 & 10'h380;
  assign T_1556 = T_1554 == 10'h0;
  assign T_1557 = Queue_1_io_deq_bits_index ^ 10'h7;
  assign T_1558 = T_1557 & 10'h380;
  assign T_1560 = T_1558 == 10'h0;
  assign T_1562 = T_1028_bits_index ^ 10'h27;
  assign T_1563 = T_1562 & 10'h380;
  assign T_1565 = T_1563 == 10'h0;
  assign T_1566 = Queue_1_io_deq_bits_index ^ 10'h27;
  assign T_1567 = T_1566 & 10'h380;
  assign T_1569 = T_1567 == 10'h0;
  assign T_1571 = T_1028_bits_index ^ 10'h42;
  assign T_1572 = T_1571 & 10'h380;
  assign T_1574 = T_1572 == 10'h0;
  assign T_1575 = Queue_1_io_deq_bits_index ^ 10'h42;
  assign T_1576 = T_1575 & 10'h380;
  assign T_1578 = T_1576 == 10'h0;
  assign T_1580 = T_1028_bits_index ^ 10'h3;
  assign T_1581 = T_1580 & 10'h380;
  assign T_1583 = T_1581 == 10'h0;
  assign T_1584 = Queue_1_io_deq_bits_index ^ 10'h3;
  assign T_1585 = T_1584 & 10'h380;
  assign T_1587 = T_1585 == 10'h0;
  assign T_1589 = T_1028_bits_index ^ 10'h50;
  assign T_1590 = T_1589 & 10'h380;
  assign T_1592 = T_1590 == 10'h0;
  assign T_1593 = Queue_1_io_deq_bits_index ^ 10'h50;
  assign T_1594 = T_1593 & 10'h380;
  assign T_1596 = T_1594 == 10'h0;
  assign T_1598 = T_1028_bits_index ^ 10'h23;
  assign T_1599 = T_1598 & 10'h380;
  assign T_1601 = T_1599 == 10'h0;
  assign T_1602 = Queue_1_io_deq_bits_index ^ 10'h23;
  assign T_1603 = T_1602 & 10'h380;
  assign T_1605 = T_1603 == 10'h0;
  assign T_1607 = T_1028_bits_index ^ 10'h12;
  assign T_1608 = T_1607 & 10'h380;
  assign T_1610 = T_1608 == 10'h0;
  assign T_1611 = Queue_1_io_deq_bits_index ^ 10'h12;
  assign T_1612 = T_1611 & 10'h380;
  assign T_1614 = T_1612 == 10'h0;
  assign T_1616 = T_1028_bits_index ^ 10'h43;
  assign T_1617 = T_1616 & 10'h380;
  assign T_1619 = T_1617 == 10'h0;
  assign T_1620 = Queue_1_io_deq_bits_index ^ 10'h43;
  assign T_1621 = T_1620 & 10'h380;
  assign T_1623 = T_1621 == 10'h0;
  assign T_1625 = T_1028_bits_index ^ 10'h10;
  assign T_1626 = T_1625 & 10'h380;
  assign T_1628 = T_1626 == 10'h0;
  assign T_1629 = Queue_1_io_deq_bits_index ^ 10'h10;
  assign T_1630 = T_1629 & 10'h380;
  assign T_1632 = T_1630 == 10'h0;
  assign T_1634 = T_1028_bits_index ^ 10'h48;
  assign T_1635 = T_1634 & 10'h380;
  assign T_1637 = T_1635 == 10'h0;
  assign T_1638 = Queue_1_io_deq_bits_index ^ 10'h48;
  assign T_1639 = T_1638 & 10'h380;
  assign T_1641 = T_1639 == 10'h0;
  assign T_1643 = T_1028_bits_index ^ 10'h2b;
  assign T_1644 = T_1643 & 10'h380;
  assign T_1646 = T_1644 == 10'h0;
  assign T_1647 = Queue_1_io_deq_bits_index ^ 10'h2b;
  assign T_1648 = T_1647 & 10'h380;
  assign T_1650 = T_1648 == 10'h0;
  assign T_1652 = T_1028_bits_index ^ 10'h28;
  assign T_1653 = T_1652 & 10'h380;
  assign T_1655 = T_1653 == 10'h0;
  assign T_1656 = Queue_1_io_deq_bits_index ^ 10'h28;
  assign T_1657 = T_1656 & 10'h380;
  assign T_1659 = T_1657 == 10'h0;
  assign T_1661 = T_1028_bits_index ^ 10'h17;
  assign T_1662 = T_1661 & 10'h380;
  assign T_1664 = T_1662 == 10'h0;
  assign T_1665 = Queue_1_io_deq_bits_index ^ 10'h17;
  assign T_1666 = T_1665 & 10'h380;
  assign T_1668 = T_1666 == 10'h0;
  assign T_1670 = T_1028_bits_index ^ 10'h8;
  assign T_1671 = T_1670 & 10'h380;
  assign T_1673 = T_1671 == 10'h0;
  assign T_1674 = Queue_1_io_deq_bits_index ^ 10'h8;
  assign T_1675 = T_1674 & 10'h380;
  assign T_1677 = T_1675 == 10'h0;
  assign T_1679 = T_1028_bits_index ^ 10'h4b;
  assign T_1680 = T_1679 & 10'h380;
  assign T_1682 = T_1680 == 10'h0;
  assign T_1683 = Queue_1_io_deq_bits_index ^ 10'h4b;
  assign T_1684 = T_1683 & 10'h380;
  assign T_1686 = T_1684 == 10'h0;
  assign T_1688 = T_1028_bits_index ^ 10'h52;
  assign T_1689 = T_1688 & 10'h380;
  assign T_1691 = T_1689 == 10'h0;
  assign T_1692 = Queue_1_io_deq_bits_index ^ 10'h52;
  assign T_1693 = T_1692 & 10'h380;
  assign T_1695 = T_1693 == 10'h0;
  assign T_1697 = T_1028_bits_index ^ 10'h24;
  assign T_1698 = T_1697 & 10'h380;
  assign T_1700 = T_1698 == 10'h0;
  assign T_1701 = Queue_1_io_deq_bits_index ^ 10'h24;
  assign T_1702 = T_1701 & 10'h380;
  assign T_1704 = T_1702 == 10'h0;
  assign T_1706 = T_1028_bits_index ^ 10'h13;
  assign T_1707 = T_1706 & 10'h380;
  assign T_1709 = T_1707 == 10'h0;
  assign T_1710 = Queue_1_io_deq_bits_index ^ 10'h13;
  assign T_1711 = T_1710 & 10'h380;
  assign T_1713 = T_1711 == 10'h0;
  assign T_1715 = T_1028_bits_index ^ 10'h4;
  assign T_1716 = T_1715 & 10'h380;
  assign T_1718 = T_1716 == 10'h0;
  assign T_1719 = Queue_1_io_deq_bits_index ^ 10'h4;
  assign T_1720 = T_1719 & 10'h380;
  assign T_1722 = T_1720 == 10'h0;
  assign T_1724 = T_1028_bits_index ^ 10'h4f;
  assign T_1725 = T_1724 & 10'h380;
  assign T_1727 = T_1725 == 10'h0;
  assign T_1728 = Queue_1_io_deq_bits_index ^ 10'h4f;
  assign T_1729 = T_1728 & 10'h380;
  assign T_1731 = T_1729 == 10'h0;
  assign T_1733 = T_1028_bits_index ^ 10'h2f;
  assign T_1734 = T_1733 & 10'h380;
  assign T_1736 = T_1734 == 10'h0;
  assign T_1737 = Queue_1_io_deq_bits_index ^ 10'h2f;
  assign T_1738 = T_1737 & 10'h380;
  assign T_1740 = T_1738 == 10'h0;
  assign T_1742 = T_1028_bits_index ^ 10'h44;
  assign T_1743 = T_1742 & 10'h380;
  assign T_1745 = T_1743 == 10'h0;
  assign T_1746 = Queue_1_io_deq_bits_index ^ 10'h44;
  assign T_1747 = T_1746 & 10'h380;
  assign T_1749 = T_1747 == 10'h0;
  assign T_1751 = T_1028_bits_index ^ 10'h53;
  assign T_1752 = T_1751 & 10'h380;
  assign T_1754 = T_1752 == 10'h0;
  assign T_1755 = Queue_1_io_deq_bits_index ^ 10'h53;
  assign T_1756 = T_1755 & 10'h380;
  assign T_1758 = T_1756 == 10'h0;
  assign T_1762_0 = T_8954;
  assign T_1762_1 = T_7574;
  assign T_1762_2 = T_8414;
  assign T_1762_3 = T_8054;
  assign T_1762_4 = T_8314;
  assign T_1762_5 = T_7974;
  assign T_1762_6 = T_8494;
  assign T_1762_7 = T_9134;
  assign T_1762_8 = T_9054;
  assign T_1762_9 = T_7694;
  assign T_1762_10 = T_8334;
  assign T_1762_11 = T_8974;
  assign T_1762_12 = T_8234;
  assign T_1762_13 = T_8874;
  assign T_1762_14 = T_9114;
  assign T_1762_15 = T_8394;
  assign T_1762_16 = T_9034;
  assign T_1762_17 = T_7614;
  assign T_1762_18 = T_8214;
  assign T_1762_19 = T_8254;
  assign T_1762_20 = T_8474;
  assign T_1762_21 = T_8854;
  assign T_1762_22 = T_8014;
  assign T_1762_23 = T_8454;
  assign T_1762_24 = T_8994;
  assign T_1762_25 = T_9194;
  assign T_1762_26 = T_9094;
  assign T_1762_27 = T_7714;
  assign T_1762_28 = T_8354;
  assign T_1762_29 = T_8894;
  assign T_1762_30 = T_7634;
  assign T_1762_31 = T_9174;
  assign T_1762_32 = T_8274;
  assign T_1762_33 = T_7934;
  assign T_1762_34 = T_8914;
  assign T_1762_35 = T_7894;
  assign T_1762_36 = T_9014;
  assign T_1762_37 = T_8434;
  assign T_1762_38 = T_8374;
  assign T_1762_39 = T_8034;
  assign T_1762_40 = T_7734;
  assign T_1762_41 = T_9074;
  assign T_1762_42 = T_9214;
  assign T_1762_43 = T_8294;
  assign T_1762_44 = T_7954;
  assign T_1762_45 = T_7654;
  assign T_1762_46 = T_9154;
  assign T_1762_47 = T_8514;
  assign T_1762_48 = T_8934;
  assign T_1762_49 = T_9234;
  assign T_1767_0 = T_8960;
  assign T_1767_1 = T_7580;
  assign T_1767_2 = T_8420;
  assign T_1767_3 = T_8060;
  assign T_1767_4 = T_8320;
  assign T_1767_5 = T_7980;
  assign T_1767_6 = T_8500;
  assign T_1767_7 = T_9140;
  assign T_1767_8 = T_9060;
  assign T_1767_9 = T_7700;
  assign T_1767_10 = T_8340;
  assign T_1767_11 = T_8980;
  assign T_1767_12 = T_8240;
  assign T_1767_13 = T_8880;
  assign T_1767_14 = T_9120;
  assign T_1767_15 = T_8400;
  assign T_1767_16 = T_9040;
  assign T_1767_17 = T_7620;
  assign T_1767_18 = T_8220;
  assign T_1767_19 = T_8260;
  assign T_1767_20 = T_8480;
  assign T_1767_21 = T_8860;
  assign T_1767_22 = T_8020;
  assign T_1767_23 = T_8460;
  assign T_1767_24 = T_9000;
  assign T_1767_25 = T_9200;
  assign T_1767_26 = T_9100;
  assign T_1767_27 = T_7720;
  assign T_1767_28 = T_8360;
  assign T_1767_29 = T_8900;
  assign T_1767_30 = T_7640;
  assign T_1767_31 = T_9180;
  assign T_1767_32 = T_8280;
  assign T_1767_33 = T_7940;
  assign T_1767_34 = T_8920;
  assign T_1767_35 = T_7900;
  assign T_1767_36 = T_9020;
  assign T_1767_37 = T_8440;
  assign T_1767_38 = T_8380;
  assign T_1767_39 = T_8040;
  assign T_1767_40 = T_7740;
  assign T_1767_41 = T_9080;
  assign T_1767_42 = T_9220;
  assign T_1767_43 = T_8300;
  assign T_1767_44 = T_7960;
  assign T_1767_45 = T_7660;
  assign T_1767_46 = T_9160;
  assign T_1767_47 = T_8520;
  assign T_1767_48 = T_8940;
  assign T_1767_49 = T_9240;
  assign T_1772_0 = 1'h1;
  assign T_1772_1 = 1'h1;
  assign T_1772_2 = 1'h1;
  assign T_1772_3 = 1'h1;
  assign T_1772_4 = 1'h1;
  assign T_1772_5 = 1'h1;
  assign T_1772_6 = 1'h1;
  assign T_1772_7 = 1'h1;
  assign T_1772_8 = 1'h1;
  assign T_1772_9 = 1'h1;
  assign T_1772_10 = 1'h1;
  assign T_1772_11 = 1'h1;
  assign T_1772_12 = 1'h1;
  assign T_1772_13 = 1'h1;
  assign T_1772_14 = 1'h1;
  assign T_1772_15 = 1'h1;
  assign T_1772_16 = 1'h1;
  assign T_1772_17 = 1'h1;
  assign T_1772_18 = 1'h1;
  assign T_1772_19 = 1'h1;
  assign T_1772_20 = 1'h1;
  assign T_1772_21 = 1'h1;
  assign T_1772_22 = 1'h1;
  assign T_1772_23 = 1'h1;
  assign T_1772_24 = 1'h1;
  assign T_1772_25 = 1'h1;
  assign T_1772_26 = 1'h1;
  assign T_1772_27 = 1'h1;
  assign T_1772_28 = 1'h1;
  assign T_1772_29 = 1'h1;
  assign T_1772_30 = 1'h1;
  assign T_1772_31 = 1'h1;
  assign T_1772_32 = 1'h1;
  assign T_1772_33 = 1'h1;
  assign T_1772_34 = 1'h1;
  assign T_1772_35 = 1'h1;
  assign T_1772_36 = 1'h1;
  assign T_1772_37 = 1'h1;
  assign T_1772_38 = 1'h1;
  assign T_1772_39 = 1'h1;
  assign T_1772_40 = 1'h1;
  assign T_1772_41 = 1'h1;
  assign T_1772_42 = 1'h1;
  assign T_1772_43 = 1'h1;
  assign T_1772_44 = 1'h1;
  assign T_1772_45 = 1'h1;
  assign T_1772_46 = 1'h1;
  assign T_1772_47 = 1'h1;
  assign T_1772_48 = 1'h1;
  assign T_1772_49 = 1'h1;
  assign T_1777_0 = 1'h1;
  assign T_1777_1 = 1'h1;
  assign T_1777_2 = 1'h1;
  assign T_1777_3 = 1'h1;
  assign T_1777_4 = 1'h1;
  assign T_1777_5 = 1'h1;
  assign T_1777_6 = 1'h1;
  assign T_1777_7 = 1'h1;
  assign T_1777_8 = 1'h1;
  assign T_1777_9 = 1'h1;
  assign T_1777_10 = 1'h1;
  assign T_1777_11 = 1'h1;
  assign T_1777_12 = 1'h1;
  assign T_1777_13 = 1'h1;
  assign T_1777_14 = 1'h1;
  assign T_1777_15 = 1'h1;
  assign T_1777_16 = 1'h1;
  assign T_1777_17 = 1'h1;
  assign T_1777_18 = 1'h1;
  assign T_1777_19 = 1'h1;
  assign T_1777_20 = 1'h1;
  assign T_1777_21 = 1'h1;
  assign T_1777_22 = 1'h1;
  assign T_1777_23 = 1'h1;
  assign T_1777_24 = 1'h1;
  assign T_1777_25 = 1'h1;
  assign T_1777_26 = 1'h1;
  assign T_1777_27 = 1'h1;
  assign T_1777_28 = 1'h1;
  assign T_1777_29 = 1'h1;
  assign T_1777_30 = 1'h1;
  assign T_1777_31 = 1'h1;
  assign T_1777_32 = 1'h1;
  assign T_1777_33 = 1'h1;
  assign T_1777_34 = 1'h1;
  assign T_1777_35 = 1'h1;
  assign T_1777_36 = 1'h1;
  assign T_1777_37 = 1'h1;
  assign T_1777_38 = 1'h1;
  assign T_1777_39 = 1'h1;
  assign T_1777_40 = 1'h1;
  assign T_1777_41 = 1'h1;
  assign T_1777_42 = 1'h1;
  assign T_1777_43 = 1'h1;
  assign T_1777_44 = 1'h1;
  assign T_1777_45 = 1'h1;
  assign T_1777_46 = 1'h1;
  assign T_1777_47 = 1'h1;
  assign T_1777_48 = 1'h1;
  assign T_1777_49 = 1'h1;
  assign T_1782_0 = 1'h1;
  assign T_1782_1 = 1'h1;
  assign T_1782_2 = 1'h1;
  assign T_1782_3 = 1'h1;
  assign T_1782_4 = 1'h1;
  assign T_1782_5 = 1'h1;
  assign T_1782_6 = 1'h1;
  assign T_1782_7 = 1'h1;
  assign T_1782_8 = 1'h1;
  assign T_1782_9 = 1'h1;
  assign T_1782_10 = 1'h1;
  assign T_1782_11 = 1'h1;
  assign T_1782_12 = 1'h1;
  assign T_1782_13 = 1'h1;
  assign T_1782_14 = 1'h1;
  assign T_1782_15 = 1'h1;
  assign T_1782_16 = 1'h1;
  assign T_1782_17 = 1'h1;
  assign T_1782_18 = 1'h1;
  assign T_1782_19 = 1'h1;
  assign T_1782_20 = 1'h1;
  assign T_1782_21 = 1'h1;
  assign T_1782_22 = 1'h1;
  assign T_1782_23 = 1'h1;
  assign T_1782_24 = 1'h1;
  assign T_1782_25 = 1'h1;
  assign T_1782_26 = 1'h1;
  assign T_1782_27 = 1'h1;
  assign T_1782_28 = 1'h1;
  assign T_1782_29 = 1'h1;
  assign T_1782_30 = 1'h1;
  assign T_1782_31 = 1'h1;
  assign T_1782_32 = 1'h1;
  assign T_1782_33 = 1'h1;
  assign T_1782_34 = 1'h1;
  assign T_1782_35 = 1'h1;
  assign T_1782_36 = 1'h1;
  assign T_1782_37 = 1'h1;
  assign T_1782_38 = 1'h1;
  assign T_1782_39 = 1'h1;
  assign T_1782_40 = 1'h1;
  assign T_1782_41 = 1'h1;
  assign T_1782_42 = 1'h1;
  assign T_1782_43 = 1'h1;
  assign T_1782_44 = 1'h1;
  assign T_1782_45 = 1'h1;
  assign T_1782_46 = 1'h1;
  assign T_1782_47 = 1'h1;
  assign T_1782_48 = 1'h1;
  assign T_1782_49 = 1'h1;
  assign T_1787_0 = 1'h1;
  assign T_1787_1 = 1'h1;
  assign T_1787_2 = 1'h1;
  assign T_1787_3 = 1'h1;
  assign T_1787_4 = 1'h1;
  assign T_1787_5 = 1'h1;
  assign T_1787_6 = 1'h1;
  assign T_1787_7 = 1'h1;
  assign T_1787_8 = 1'h1;
  assign T_1787_9 = 1'h1;
  assign T_1787_10 = 1'h1;
  assign T_1787_11 = 1'h1;
  assign T_1787_12 = 1'h1;
  assign T_1787_13 = 1'h1;
  assign T_1787_14 = 1'h1;
  assign T_1787_15 = 1'h1;
  assign T_1787_16 = 1'h1;
  assign T_1787_17 = 1'h1;
  assign T_1787_18 = 1'h1;
  assign T_1787_19 = 1'h1;
  assign T_1787_20 = 1'h1;
  assign T_1787_21 = 1'h1;
  assign T_1787_22 = 1'h1;
  assign T_1787_23 = 1'h1;
  assign T_1787_24 = 1'h1;
  assign T_1787_25 = 1'h1;
  assign T_1787_26 = 1'h1;
  assign T_1787_27 = 1'h1;
  assign T_1787_28 = 1'h1;
  assign T_1787_29 = 1'h1;
  assign T_1787_30 = 1'h1;
  assign T_1787_31 = 1'h1;
  assign T_1787_32 = 1'h1;
  assign T_1787_33 = 1'h1;
  assign T_1787_34 = 1'h1;
  assign T_1787_35 = 1'h1;
  assign T_1787_36 = 1'h1;
  assign T_1787_37 = 1'h1;
  assign T_1787_38 = 1'h1;
  assign T_1787_39 = 1'h1;
  assign T_1787_40 = 1'h1;
  assign T_1787_41 = 1'h1;
  assign T_1787_42 = 1'h1;
  assign T_1787_43 = 1'h1;
  assign T_1787_44 = 1'h1;
  assign T_1787_45 = 1'h1;
  assign T_1787_46 = 1'h1;
  assign T_1787_47 = 1'h1;
  assign T_1787_48 = 1'h1;
  assign T_1787_49 = 1'h1;
  assign T_1792_0 = T_8964;
  assign T_1792_1 = T_7584;
  assign T_1792_2 = T_8424;
  assign T_1792_3 = T_8064;
  assign T_1792_4 = T_8324;
  assign T_1792_5 = T_7984;
  assign T_1792_6 = T_8504;
  assign T_1792_7 = T_9144;
  assign T_1792_8 = T_9064;
  assign T_1792_9 = T_7704;
  assign T_1792_10 = T_8344;
  assign T_1792_11 = T_8984;
  assign T_1792_12 = T_8244;
  assign T_1792_13 = T_8884;
  assign T_1792_14 = T_9124;
  assign T_1792_15 = T_8404;
  assign T_1792_16 = T_9044;
  assign T_1792_17 = T_7624;
  assign T_1792_18 = T_8224;
  assign T_1792_19 = T_8264;
  assign T_1792_20 = T_8484;
  assign T_1792_21 = T_8864;
  assign T_1792_22 = T_8024;
  assign T_1792_23 = T_8464;
  assign T_1792_24 = T_9004;
  assign T_1792_25 = T_9204;
  assign T_1792_26 = T_9104;
  assign T_1792_27 = T_7724;
  assign T_1792_28 = T_8364;
  assign T_1792_29 = T_8904;
  assign T_1792_30 = T_7644;
  assign T_1792_31 = T_9184;
  assign T_1792_32 = T_8284;
  assign T_1792_33 = T_7944;
  assign T_1792_34 = T_8924;
  assign T_1792_35 = T_7904;
  assign T_1792_36 = T_9024;
  assign T_1792_37 = T_8444;
  assign T_1792_38 = T_8384;
  assign T_1792_39 = T_8044;
  assign T_1792_40 = T_7744;
  assign T_1792_41 = T_9084;
  assign T_1792_42 = T_9224;
  assign T_1792_43 = T_8304;
  assign T_1792_44 = T_7964;
  assign T_1792_45 = T_7664;
  assign T_1792_46 = T_9164;
  assign T_1792_47 = T_8524;
  assign T_1792_48 = T_8944;
  assign T_1792_49 = T_9244;
  assign T_1797_0 = T_8970;
  assign T_1797_1 = T_7590;
  assign T_1797_2 = T_8430;
  assign T_1797_3 = T_8070;
  assign T_1797_4 = T_8330;
  assign T_1797_5 = T_7990;
  assign T_1797_6 = T_8510;
  assign T_1797_7 = T_9150;
  assign T_1797_8 = T_9070;
  assign T_1797_9 = T_7710;
  assign T_1797_10 = T_8350;
  assign T_1797_11 = T_8990;
  assign T_1797_12 = T_8250;
  assign T_1797_13 = T_8890;
  assign T_1797_14 = T_9130;
  assign T_1797_15 = T_8410;
  assign T_1797_16 = T_9050;
  assign T_1797_17 = T_7630;
  assign T_1797_18 = T_8230;
  assign T_1797_19 = T_8270;
  assign T_1797_20 = T_8490;
  assign T_1797_21 = T_8870;
  assign T_1797_22 = T_8030;
  assign T_1797_23 = T_8470;
  assign T_1797_24 = T_9010;
  assign T_1797_25 = T_9210;
  assign T_1797_26 = T_9110;
  assign T_1797_27 = T_7730;
  assign T_1797_28 = T_8370;
  assign T_1797_29 = T_8910;
  assign T_1797_30 = T_7650;
  assign T_1797_31 = T_9190;
  assign T_1797_32 = T_8290;
  assign T_1797_33 = T_7950;
  assign T_1797_34 = T_8930;
  assign T_1797_35 = T_7910;
  assign T_1797_36 = T_9030;
  assign T_1797_37 = T_8450;
  assign T_1797_38 = T_8390;
  assign T_1797_39 = T_8050;
  assign T_1797_40 = T_7750;
  assign T_1797_41 = T_9090;
  assign T_1797_42 = T_9230;
  assign T_1797_43 = T_8310;
  assign T_1797_44 = T_7970;
  assign T_1797_45 = T_7670;
  assign T_1797_46 = T_9170;
  assign T_1797_47 = T_8530;
  assign T_1797_48 = T_8950;
  assign T_1797_49 = T_9250;
  assign T_2462 = Queue_1_io_deq_bits_mask[0];
  assign T_2463 = Queue_1_io_deq_bits_mask[1];
  assign T_2464 = Queue_1_io_deq_bits_mask[2];
  assign T_2465 = Queue_1_io_deq_bits_mask[3];
  assign T_2469 = T_2462 ? 8'hff : 8'h0;
  assign T_2473 = T_2463 ? 8'hff : 8'h0;
  assign T_2477 = T_2464 ? 8'hff : 8'h0;
  assign T_2481 = T_2465 ? 8'hff : 8'h0;
  assign T_2482 = {T_2473,T_2469};
  assign T_2483 = {T_2481,T_2477};
  assign T_2484 = {T_2483,T_2482};
  assign T_2496 = ~ T_2484;
  assign T_2498 = T_2496 == 32'h0;
  assign T_2504 = T_1797_0 & T_2498;
  assign T_2505 = Queue_1_io_deq_bits_data;
  assign T_2520 = pmu_io_regs_wakeupProgram_5_read;
  assign T_2544 = T_1797_1 & T_2498;
  assign T_2560 = wdog_io_regs_cfg_read;
  assign T_2584 = T_1797_2 & T_2498;
  assign GEN_6 = T_2584 ? T_2505 : backupRegs_10;
  assign T_2624 = T_1797_3 & T_2498;
  assign T_2640 = rtc_io_regs_cmp_0_read;
  assign T_2664 = T_1797_4 & T_2498;
  assign GEN_7 = T_2664 ? T_2505 : backupRegs_5;
  assign T_2704 = T_1797_5 & T_2498;
  assign T_2720 = rtc_io_regs_s_read;
  assign T_2744 = T_1797_6 & T_2498;
  assign GEN_8 = T_2744 ? T_2505 : backupRegs_14;
  assign T_2784 = T_1797_7 & T_2498;
  assign T_2800 = pmu_io_regs_sleepProgram_6_read;
  assign T_2824 = T_1797_8 & T_2498;
  assign T_2840 = pmu_io_regs_sleepProgram_2_read;
  assign T_2864 = T_1797_9 & T_2498;
  assign T_2880 = wdog_io_regs_feed_read;
  assign T_2904 = T_1797_10 & T_2498;
  assign GEN_9 = T_2904 ? T_2505 : backupRegs_6;
  assign T_2944 = T_1797_11 & T_2498;
  assign T_2960 = pmu_io_regs_wakeupProgram_6_read;
  assign T_2984 = T_1797_12 & T_2498;
  assign GEN_10 = T_2984 ? T_2505 : backupRegs_1;
  assign T_3024 = T_1797_13 & T_2498;
  assign T_3040 = pmu_io_regs_wakeupProgram_1_read;
  assign T_3064 = T_1797_14 & T_2498;
  assign T_3080 = pmu_io_regs_sleepProgram_5_read;
  assign T_3104 = T_1797_15 & T_2498;
  assign GEN_11 = T_3104 ? T_2505 : backupRegs_9;
  assign T_3144 = T_1797_16 & T_2498;
  assign T_3160 = pmu_io_regs_sleepProgram_1_read;
  assign T_3184 = T_1797_17 & T_2498;
  assign T_3200 = wdog_io_regs_countLo_read;
  assign T_3224 = T_1797_18 & T_2498;
  assign GEN_12 = T_3224 ? T_2505 : backupRegs_0;
  assign T_3264 = T_1797_19 & T_2498;
  assign GEN_13 = T_3264 ? T_2505 : backupRegs_2;
  assign T_3304 = T_1797_20 & T_2498;
  assign GEN_14 = T_3304 ? T_2505 : backupRegs_13;
  assign T_3344 = T_1797_21 & T_2498;
  assign T_3360 = pmu_io_regs_wakeupProgram_0_read;
  assign T_3384 = T_1797_22 & T_2498;
  assign T_3400 = rtc_io_regs_feed_read;
  assign T_3424 = T_1797_23 & T_2498;
  assign GEN_15 = T_3424 ? T_2505 : backupRegs_12;
  assign T_3464 = T_1797_24 & T_2498;
  assign T_3480 = pmu_io_regs_wakeupProgram_7_read;
  assign T_3504 = T_1797_25 & T_2498;
  assign T_3520 = pmu_io_regs_cause_read;
  assign T_3544 = T_1797_26 & T_2498;
  assign T_3560 = pmu_io_regs_sleepProgram_4_read;
  assign T_3584 = T_1797_27 & T_2498;
  assign T_3600 = wdog_io_regs_key_read;
  assign T_3624 = T_1797_28 & T_2498;
  assign GEN_16 = T_3624 ? T_2505 : backupRegs_7;
  assign T_3664 = T_1797_29 & T_2498;
  assign T_3680 = pmu_io_regs_wakeupProgram_2_read;
  assign T_3704 = T_1797_30 & T_2498;
  assign T_3720 = wdog_io_regs_countHi_read;
  assign T_3732 = T_2484[3:0];
  assign T_3736 = ~ T_3732;
  assign T_3738 = T_3736 == 4'h0;
  assign T_3744 = T_1797_31 & T_3738;
  assign T_3745 = Queue_1_io_deq_bits_data[3:0];
  assign T_3760 = pmu_io_regs_ie_read;
  assign T_3784 = T_1797_32 & T_2498;
  assign GEN_17 = T_3784 ? T_2505 : backupRegs_3;
  assign T_3824 = T_1797_33 & T_2498;
  assign T_3840 = rtc_io_regs_countLo_read;
  assign T_3864 = T_1797_34 & T_2498;
  assign T_3880 = pmu_io_regs_wakeupProgram_3_read;
  assign T_3904 = T_1797_35 & T_2498;
  assign T_3920 = rtc_io_regs_cfg_read;
  assign T_3944 = T_1797_36 & T_2498;
  assign T_3960 = pmu_io_regs_sleepProgram_0_read;
  assign T_3984 = T_1797_37 & T_2498;
  assign GEN_18 = T_3984 ? T_2505 : backupRegs_11;
  assign T_4024 = T_1797_38 & T_2498;
  assign GEN_19 = T_4024 ? T_2505 : backupRegs_8;
  assign T_4064 = T_1797_39 & T_2498;
  assign T_4080 = rtc_io_regs_key_read;
  assign T_4092 = T_2484[15:0];
  assign T_4096 = ~ T_4092;
  assign T_4098 = T_4096 == 16'h0;
  assign T_4104 = T_1797_40 & T_4098;
  assign T_4105 = Queue_1_io_deq_bits_data[15:0];
  assign T_4120 = wdog_io_regs_cmp_0_read;
  assign T_4144 = T_1797_41 & T_2498;
  assign T_4160 = pmu_io_regs_sleepProgram_3_read;
  assign T_4184 = T_1797_42 & T_2498;
  assign T_4200 = pmu_io_regs_sleep_read;
  assign T_4224 = T_1797_43 & T_2498;
  assign GEN_20 = T_4224 ? T_2505 : backupRegs_4;
  assign T_4264 = T_1797_44 & T_2498;
  assign T_4280 = rtc_io_regs_countHi_read;
  assign T_4304 = T_1797_45 & T_4098;
  assign T_4320 = wdog_io_regs_s_read;
  assign T_4344 = T_1797_46 & T_2498;
  assign T_4360 = pmu_io_regs_sleepProgram_7_read;
  assign T_4384 = T_1797_47 & T_2498;
  assign GEN_21 = T_4384 ? T_2505 : backupRegs_15;
  assign T_4424 = T_1797_48 & T_2498;
  assign T_4440 = pmu_io_regs_wakeupProgram_4_read;
  assign T_4464 = T_1797_49 & T_2498;
  assign T_4480 = pmu_io_regs_key_read;
  assign T_4486 = T_1322 == 1'h0;
  assign T_4488 = T_4486 | T_1772_1;
  assign T_4493 = T_1466 == 1'h0;
  assign T_4495 = T_4493 | T_1772_17;
  assign T_4497 = T_1583 == 1'h0;
  assign T_4499 = T_4497 | T_1772_30;
  assign T_4501 = T_1718 == 1'h0;
  assign T_4503 = T_4501 | T_1772_45;
  assign T_4508 = T_1394 == 1'h0;
  assign T_4510 = T_4508 | T_1772_9;
  assign T_4512 = T_1556 == 1'h0;
  assign T_4514 = T_4512 | T_1772_27;
  assign T_4516 = T_1673 == 1'h0;
  assign T_4518 = T_4516 | T_1772_40;
  assign T_4541 = T_1628 == 1'h0;
  assign T_4543 = T_4541 | T_1772_35;
  assign T_4548 = T_1610 == 1'h0;
  assign T_4550 = T_4548 | T_1772_33;
  assign T_4552 = T_1709 == 1'h0;
  assign T_4554 = T_4552 | T_1772_44;
  assign T_4556 = T_1358 == 1'h0;
  assign T_4558 = T_4556 | T_1772_5;
  assign T_4563 = T_1511 == 1'h0;
  assign T_4565 = T_4563 | T_1772_22;
  assign T_4567 = T_1664 == 1'h0;
  assign T_4569 = T_4567 | T_1772_39;
  assign T_4571 = T_1340 == 1'h0;
  assign T_4573 = T_4571 | T_1772_3;
  assign T_4596 = T_1475 == 1'h0;
  assign T_4598 = T_4596 | T_1772_18;
  assign T_4600 = T_1421 == 1'h0;
  assign T_4602 = T_4600 | T_1772_12;
  assign T_4604 = T_1484 == 1'h0;
  assign T_4606 = T_4604 | T_1772_19;
  assign T_4608 = T_1601 == 1'h0;
  assign T_4610 = T_4608 | T_1772_32;
  assign T_4612 = T_1700 == 1'h0;
  assign T_4614 = T_4612 | T_1772_43;
  assign T_4616 = T_1349 == 1'h0;
  assign T_4618 = T_4616 | T_1772_4;
  assign T_4620 = T_1403 == 1'h0;
  assign T_4622 = T_4620 | T_1772_10;
  assign T_4624 = T_1565 == 1'h0;
  assign T_4626 = T_4624 | T_1772_28;
  assign T_4628 = T_1655 == 1'h0;
  assign T_4630 = T_4628 | T_1772_38;
  assign T_4632 = T_1448 == 1'h0;
  assign T_4634 = T_4632 | T_1772_15;
  assign T_4636 = T_1331 == 1'h0;
  assign T_4638 = T_4636 | T_1772_2;
  assign T_4640 = T_1646 == 1'h0;
  assign T_4642 = T_4640 | T_1772_37;
  assign T_4644 = T_1520 == 1'h0;
  assign T_4646 = T_4644 | T_1772_23;
  assign T_4648 = T_1493 == 1'h0;
  assign T_4650 = T_4648 | T_1772_20;
  assign T_4652 = T_1367 == 1'h0;
  assign T_4654 = T_4652 | T_1772_6;
  assign T_4656 = T_1736 == 1'h0;
  assign T_4658 = T_4656 | T_1772_47;
  assign T_4708 = T_1502 == 1'h0;
  assign T_4710 = T_4708 | T_1772_21;
  assign T_4712 = T_1430 == 1'h0;
  assign T_4714 = T_4712 | T_1772_13;
  assign T_4716 = T_1574 == 1'h0;
  assign T_4718 = T_4716 | T_1772_29;
  assign T_4720 = T_1619 == 1'h0;
  assign T_4722 = T_4720 | T_1772_34;
  assign T_4724 = T_1745 == 1'h0;
  assign T_4726 = T_4724 | T_1772_48;
  assign T_4728 = T_1313 == 1'h0;
  assign T_4730 = T_4728 | T_1772_0;
  assign T_4732 = T_1412 == 1'h0;
  assign T_4734 = T_4732 | T_1772_11;
  assign T_4736 = T_1529 == 1'h0;
  assign T_4738 = T_4736 | T_1772_24;
  assign T_4740 = T_1637 == 1'h0;
  assign T_4742 = T_4740 | T_1772_36;
  assign T_4744 = T_1457 == 1'h0;
  assign T_4746 = T_4744 | T_1772_16;
  assign T_4748 = T_1385 == 1'h0;
  assign T_4750 = T_4748 | T_1772_8;
  assign T_4752 = T_1682 == 1'h0;
  assign T_4754 = T_4752 | T_1772_41;
  assign T_4756 = T_1547 == 1'h0;
  assign T_4758 = T_4756 | T_1772_26;
  assign T_4760 = T_1439 == 1'h0;
  assign T_4762 = T_4760 | T_1772_14;
  assign T_4764 = T_1376 == 1'h0;
  assign T_4766 = T_4764 | T_1772_7;
  assign T_4768 = T_1727 == 1'h0;
  assign T_4770 = T_4768 | T_1772_46;
  assign T_4772 = T_1592 == 1'h0;
  assign T_4774 = T_4772 | T_1772_31;
  assign T_4776 = T_1538 == 1'h0;
  assign T_4778 = T_4776 | T_1772_25;
  assign T_4780 = T_1691 == 1'h0;
  assign T_4782 = T_4780 | T_1772_42;
  assign T_4784 = T_1754 == 1'h0;
  assign T_4786 = T_4784 | T_1772_49;
  assign T_5050_0 = T_4488;
  assign T_5050_1 = 1'h1;
  assign T_5050_2 = T_4495;
  assign T_5050_3 = T_4499;
  assign T_5050_4 = T_4503;
  assign T_5050_5 = 1'h1;
  assign T_5050_6 = T_4510;
  assign T_5050_7 = T_4514;
  assign T_5050_8 = T_4518;
  assign T_5050_9 = 1'h1;
  assign T_5050_10 = 1'h1;
  assign T_5050_11 = 1'h1;
  assign T_5050_12 = 1'h1;
  assign T_5050_13 = 1'h1;
  assign T_5050_14 = 1'h1;
  assign T_5050_15 = 1'h1;
  assign T_5050_16 = T_4543;
  assign T_5050_17 = 1'h1;
  assign T_5050_18 = T_4550;
  assign T_5050_19 = T_4554;
  assign T_5050_20 = T_4558;
  assign T_5050_21 = 1'h1;
  assign T_5050_22 = T_4565;
  assign T_5050_23 = T_4569;
  assign T_5050_24 = T_4573;
  assign T_5050_25 = 1'h1;
  assign T_5050_26 = 1'h1;
  assign T_5050_27 = 1'h1;
  assign T_5050_28 = 1'h1;
  assign T_5050_29 = 1'h1;
  assign T_5050_30 = 1'h1;
  assign T_5050_31 = 1'h1;
  assign T_5050_32 = T_4598;
  assign T_5050_33 = T_4602;
  assign T_5050_34 = T_4606;
  assign T_5050_35 = T_4610;
  assign T_5050_36 = T_4614;
  assign T_5050_37 = T_4618;
  assign T_5050_38 = T_4622;
  assign T_5050_39 = T_4626;
  assign T_5050_40 = T_4630;
  assign T_5050_41 = T_4634;
  assign T_5050_42 = T_4638;
  assign T_5050_43 = T_4642;
  assign T_5050_44 = T_4646;
  assign T_5050_45 = T_4650;
  assign T_5050_46 = T_4654;
  assign T_5050_47 = T_4658;
  assign T_5050_48 = 1'h1;
  assign T_5050_49 = 1'h1;
  assign T_5050_50 = 1'h1;
  assign T_5050_51 = 1'h1;
  assign T_5050_52 = 1'h1;
  assign T_5050_53 = 1'h1;
  assign T_5050_54 = 1'h1;
  assign T_5050_55 = 1'h1;
  assign T_5050_56 = 1'h1;
  assign T_5050_57 = 1'h1;
  assign T_5050_58 = 1'h1;
  assign T_5050_59 = 1'h1;
  assign T_5050_60 = 1'h1;
  assign T_5050_61 = 1'h1;
  assign T_5050_62 = 1'h1;
  assign T_5050_63 = 1'h1;
  assign T_5050_64 = T_4710;
  assign T_5050_65 = T_4714;
  assign T_5050_66 = T_4718;
  assign T_5050_67 = T_4722;
  assign T_5050_68 = T_4726;
  assign T_5050_69 = T_4730;
  assign T_5050_70 = T_4734;
  assign T_5050_71 = T_4738;
  assign T_5050_72 = T_4742;
  assign T_5050_73 = T_4746;
  assign T_5050_74 = T_4750;
  assign T_5050_75 = T_4754;
  assign T_5050_76 = T_4758;
  assign T_5050_77 = T_4762;
  assign T_5050_78 = T_4766;
  assign T_5050_79 = T_4770;
  assign T_5050_80 = T_4774;
  assign T_5050_81 = T_4778;
  assign T_5050_82 = T_4782;
  assign T_5050_83 = T_4786;
  assign T_5050_84 = 1'h1;
  assign T_5050_85 = 1'h1;
  assign T_5050_86 = 1'h1;
  assign T_5050_87 = 1'h1;
  assign T_5050_88 = 1'h1;
  assign T_5050_89 = 1'h1;
  assign T_5050_90 = 1'h1;
  assign T_5050_91 = 1'h1;
  assign T_5050_92 = 1'h1;
  assign T_5050_93 = 1'h1;
  assign T_5050_94 = 1'h1;
  assign T_5050_95 = 1'h1;
  assign T_5050_96 = 1'h1;
  assign T_5050_97 = 1'h1;
  assign T_5050_98 = 1'h1;
  assign T_5050_99 = 1'h1;
  assign T_5050_100 = 1'h1;
  assign T_5050_101 = 1'h1;
  assign T_5050_102 = 1'h1;
  assign T_5050_103 = 1'h1;
  assign T_5050_104 = 1'h1;
  assign T_5050_105 = 1'h1;
  assign T_5050_106 = 1'h1;
  assign T_5050_107 = 1'h1;
  assign T_5050_108 = 1'h1;
  assign T_5050_109 = 1'h1;
  assign T_5050_110 = 1'h1;
  assign T_5050_111 = 1'h1;
  assign T_5050_112 = 1'h1;
  assign T_5050_113 = 1'h1;
  assign T_5050_114 = 1'h1;
  assign T_5050_115 = 1'h1;
  assign T_5050_116 = 1'h1;
  assign T_5050_117 = 1'h1;
  assign T_5050_118 = 1'h1;
  assign T_5050_119 = 1'h1;
  assign T_5050_120 = 1'h1;
  assign T_5050_121 = 1'h1;
  assign T_5050_122 = 1'h1;
  assign T_5050_123 = 1'h1;
  assign T_5050_124 = 1'h1;
  assign T_5050_125 = 1'h1;
  assign T_5050_126 = 1'h1;
  assign T_5050_127 = 1'h1;
  assign T_5184 = T_4486 | T_1777_1;
  assign T_5191 = T_4493 | T_1777_17;
  assign T_5195 = T_4497 | T_1777_30;
  assign T_5199 = T_4501 | T_1777_45;
  assign T_5206 = T_4508 | T_1777_9;
  assign T_5210 = T_4512 | T_1777_27;
  assign T_5214 = T_4516 | T_1777_40;
  assign T_5239 = T_4541 | T_1777_35;
  assign T_5246 = T_4548 | T_1777_33;
  assign T_5250 = T_4552 | T_1777_44;
  assign T_5254 = T_4556 | T_1777_5;
  assign T_5261 = T_4563 | T_1777_22;
  assign T_5265 = T_4567 | T_1777_39;
  assign T_5269 = T_4571 | T_1777_3;
  assign T_5294 = T_4596 | T_1777_18;
  assign T_5298 = T_4600 | T_1777_12;
  assign T_5302 = T_4604 | T_1777_19;
  assign T_5306 = T_4608 | T_1777_32;
  assign T_5310 = T_4612 | T_1777_43;
  assign T_5314 = T_4616 | T_1777_4;
  assign T_5318 = T_4620 | T_1777_10;
  assign T_5322 = T_4624 | T_1777_28;
  assign T_5326 = T_4628 | T_1777_38;
  assign T_5330 = T_4632 | T_1777_15;
  assign T_5334 = T_4636 | T_1777_2;
  assign T_5338 = T_4640 | T_1777_37;
  assign T_5342 = T_4644 | T_1777_23;
  assign T_5346 = T_4648 | T_1777_20;
  assign T_5350 = T_4652 | T_1777_6;
  assign T_5354 = T_4656 | T_1777_47;
  assign T_5406 = T_4708 | T_1777_21;
  assign T_5410 = T_4712 | T_1777_13;
  assign T_5414 = T_4716 | T_1777_29;
  assign T_5418 = T_4720 | T_1777_34;
  assign T_5422 = T_4724 | T_1777_48;
  assign T_5426 = T_4728 | T_1777_0;
  assign T_5430 = T_4732 | T_1777_11;
  assign T_5434 = T_4736 | T_1777_24;
  assign T_5438 = T_4740 | T_1777_36;
  assign T_5442 = T_4744 | T_1777_16;
  assign T_5446 = T_4748 | T_1777_8;
  assign T_5450 = T_4752 | T_1777_41;
  assign T_5454 = T_4756 | T_1777_26;
  assign T_5458 = T_4760 | T_1777_14;
  assign T_5462 = T_4764 | T_1777_7;
  assign T_5466 = T_4768 | T_1777_46;
  assign T_5470 = T_4772 | T_1777_31;
  assign T_5474 = T_4776 | T_1777_25;
  assign T_5478 = T_4780 | T_1777_42;
  assign T_5482 = T_4784 | T_1777_49;
  assign T_5746_0 = T_5184;
  assign T_5746_1 = 1'h1;
  assign T_5746_2 = T_5191;
  assign T_5746_3 = T_5195;
  assign T_5746_4 = T_5199;
  assign T_5746_5 = 1'h1;
  assign T_5746_6 = T_5206;
  assign T_5746_7 = T_5210;
  assign T_5746_8 = T_5214;
  assign T_5746_9 = 1'h1;
  assign T_5746_10 = 1'h1;
  assign T_5746_11 = 1'h1;
  assign T_5746_12 = 1'h1;
  assign T_5746_13 = 1'h1;
  assign T_5746_14 = 1'h1;
  assign T_5746_15 = 1'h1;
  assign T_5746_16 = T_5239;
  assign T_5746_17 = 1'h1;
  assign T_5746_18 = T_5246;
  assign T_5746_19 = T_5250;
  assign T_5746_20 = T_5254;
  assign T_5746_21 = 1'h1;
  assign T_5746_22 = T_5261;
  assign T_5746_23 = T_5265;
  assign T_5746_24 = T_5269;
  assign T_5746_25 = 1'h1;
  assign T_5746_26 = 1'h1;
  assign T_5746_27 = 1'h1;
  assign T_5746_28 = 1'h1;
  assign T_5746_29 = 1'h1;
  assign T_5746_30 = 1'h1;
  assign T_5746_31 = 1'h1;
  assign T_5746_32 = T_5294;
  assign T_5746_33 = T_5298;
  assign T_5746_34 = T_5302;
  assign T_5746_35 = T_5306;
  assign T_5746_36 = T_5310;
  assign T_5746_37 = T_5314;
  assign T_5746_38 = T_5318;
  assign T_5746_39 = T_5322;
  assign T_5746_40 = T_5326;
  assign T_5746_41 = T_5330;
  assign T_5746_42 = T_5334;
  assign T_5746_43 = T_5338;
  assign T_5746_44 = T_5342;
  assign T_5746_45 = T_5346;
  assign T_5746_46 = T_5350;
  assign T_5746_47 = T_5354;
  assign T_5746_48 = 1'h1;
  assign T_5746_49 = 1'h1;
  assign T_5746_50 = 1'h1;
  assign T_5746_51 = 1'h1;
  assign T_5746_52 = 1'h1;
  assign T_5746_53 = 1'h1;
  assign T_5746_54 = 1'h1;
  assign T_5746_55 = 1'h1;
  assign T_5746_56 = 1'h1;
  assign T_5746_57 = 1'h1;
  assign T_5746_58 = 1'h1;
  assign T_5746_59 = 1'h1;
  assign T_5746_60 = 1'h1;
  assign T_5746_61 = 1'h1;
  assign T_5746_62 = 1'h1;
  assign T_5746_63 = 1'h1;
  assign T_5746_64 = T_5406;
  assign T_5746_65 = T_5410;
  assign T_5746_66 = T_5414;
  assign T_5746_67 = T_5418;
  assign T_5746_68 = T_5422;
  assign T_5746_69 = T_5426;
  assign T_5746_70 = T_5430;
  assign T_5746_71 = T_5434;
  assign T_5746_72 = T_5438;
  assign T_5746_73 = T_5442;
  assign T_5746_74 = T_5446;
  assign T_5746_75 = T_5450;
  assign T_5746_76 = T_5454;
  assign T_5746_77 = T_5458;
  assign T_5746_78 = T_5462;
  assign T_5746_79 = T_5466;
  assign T_5746_80 = T_5470;
  assign T_5746_81 = T_5474;
  assign T_5746_82 = T_5478;
  assign T_5746_83 = T_5482;
  assign T_5746_84 = 1'h1;
  assign T_5746_85 = 1'h1;
  assign T_5746_86 = 1'h1;
  assign T_5746_87 = 1'h1;
  assign T_5746_88 = 1'h1;
  assign T_5746_89 = 1'h1;
  assign T_5746_90 = 1'h1;
  assign T_5746_91 = 1'h1;
  assign T_5746_92 = 1'h1;
  assign T_5746_93 = 1'h1;
  assign T_5746_94 = 1'h1;
  assign T_5746_95 = 1'h1;
  assign T_5746_96 = 1'h1;
  assign T_5746_97 = 1'h1;
  assign T_5746_98 = 1'h1;
  assign T_5746_99 = 1'h1;
  assign T_5746_100 = 1'h1;
  assign T_5746_101 = 1'h1;
  assign T_5746_102 = 1'h1;
  assign T_5746_103 = 1'h1;
  assign T_5746_104 = 1'h1;
  assign T_5746_105 = 1'h1;
  assign T_5746_106 = 1'h1;
  assign T_5746_107 = 1'h1;
  assign T_5746_108 = 1'h1;
  assign T_5746_109 = 1'h1;
  assign T_5746_110 = 1'h1;
  assign T_5746_111 = 1'h1;
  assign T_5746_112 = 1'h1;
  assign T_5746_113 = 1'h1;
  assign T_5746_114 = 1'h1;
  assign T_5746_115 = 1'h1;
  assign T_5746_116 = 1'h1;
  assign T_5746_117 = 1'h1;
  assign T_5746_118 = 1'h1;
  assign T_5746_119 = 1'h1;
  assign T_5746_120 = 1'h1;
  assign T_5746_121 = 1'h1;
  assign T_5746_122 = 1'h1;
  assign T_5746_123 = 1'h1;
  assign T_5746_124 = 1'h1;
  assign T_5746_125 = 1'h1;
  assign T_5746_126 = 1'h1;
  assign T_5746_127 = 1'h1;
  assign T_5878 = T_1326 == 1'h0;
  assign T_5880 = T_5878 | T_1782_1;
  assign T_5885 = T_1470 == 1'h0;
  assign T_5887 = T_5885 | T_1782_17;
  assign T_5889 = T_1587 == 1'h0;
  assign T_5891 = T_5889 | T_1782_30;
  assign T_5893 = T_1722 == 1'h0;
  assign T_5895 = T_5893 | T_1782_45;
  assign T_5900 = T_1398 == 1'h0;
  assign T_5902 = T_5900 | T_1782_9;
  assign T_5904 = T_1560 == 1'h0;
  assign T_5906 = T_5904 | T_1782_27;
  assign T_5908 = T_1677 == 1'h0;
  assign T_5910 = T_5908 | T_1782_40;
  assign T_5933 = T_1632 == 1'h0;
  assign T_5935 = T_5933 | T_1782_35;
  assign T_5940 = T_1614 == 1'h0;
  assign T_5942 = T_5940 | T_1782_33;
  assign T_5944 = T_1713 == 1'h0;
  assign T_5946 = T_5944 | T_1782_44;
  assign T_5948 = T_1362 == 1'h0;
  assign T_5950 = T_5948 | T_1782_5;
  assign T_5955 = T_1515 == 1'h0;
  assign T_5957 = T_5955 | T_1782_22;
  assign T_5959 = T_1668 == 1'h0;
  assign T_5961 = T_5959 | T_1782_39;
  assign T_5963 = T_1344 == 1'h0;
  assign T_5965 = T_5963 | T_1782_3;
  assign T_5988 = T_1479 == 1'h0;
  assign T_5990 = T_5988 | T_1782_18;
  assign T_5992 = T_1425 == 1'h0;
  assign T_5994 = T_5992 | T_1782_12;
  assign T_5996 = T_1488 == 1'h0;
  assign T_5998 = T_5996 | T_1782_19;
  assign T_6000 = T_1605 == 1'h0;
  assign T_6002 = T_6000 | T_1782_32;
  assign T_6004 = T_1704 == 1'h0;
  assign T_6006 = T_6004 | T_1782_43;
  assign T_6008 = T_1353 == 1'h0;
  assign T_6010 = T_6008 | T_1782_4;
  assign T_6012 = T_1407 == 1'h0;
  assign T_6014 = T_6012 | T_1782_10;
  assign T_6016 = T_1569 == 1'h0;
  assign T_6018 = T_6016 | T_1782_28;
  assign T_6020 = T_1659 == 1'h0;
  assign T_6022 = T_6020 | T_1782_38;
  assign T_6024 = T_1452 == 1'h0;
  assign T_6026 = T_6024 | T_1782_15;
  assign T_6028 = T_1335 == 1'h0;
  assign T_6030 = T_6028 | T_1782_2;
  assign T_6032 = T_1650 == 1'h0;
  assign T_6034 = T_6032 | T_1782_37;
  assign T_6036 = T_1524 == 1'h0;
  assign T_6038 = T_6036 | T_1782_23;
  assign T_6040 = T_1497 == 1'h0;
  assign T_6042 = T_6040 | T_1782_20;
  assign T_6044 = T_1371 == 1'h0;
  assign T_6046 = T_6044 | T_1782_6;
  assign T_6048 = T_1740 == 1'h0;
  assign T_6050 = T_6048 | T_1782_47;
  assign T_6100 = T_1506 == 1'h0;
  assign T_6102 = T_6100 | T_1782_21;
  assign T_6104 = T_1434 == 1'h0;
  assign T_6106 = T_6104 | T_1782_13;
  assign T_6108 = T_1578 == 1'h0;
  assign T_6110 = T_6108 | T_1782_29;
  assign T_6112 = T_1623 == 1'h0;
  assign T_6114 = T_6112 | T_1782_34;
  assign T_6116 = T_1749 == 1'h0;
  assign T_6118 = T_6116 | T_1782_48;
  assign T_6120 = T_1317 == 1'h0;
  assign T_6122 = T_6120 | T_1782_0;
  assign T_6124 = T_1416 == 1'h0;
  assign T_6126 = T_6124 | T_1782_11;
  assign T_6128 = T_1533 == 1'h0;
  assign T_6130 = T_6128 | T_1782_24;
  assign T_6132 = T_1641 == 1'h0;
  assign T_6134 = T_6132 | T_1782_36;
  assign T_6136 = T_1461 == 1'h0;
  assign T_6138 = T_6136 | T_1782_16;
  assign T_6140 = T_1389 == 1'h0;
  assign T_6142 = T_6140 | T_1782_8;
  assign T_6144 = T_1686 == 1'h0;
  assign T_6146 = T_6144 | T_1782_41;
  assign T_6148 = T_1551 == 1'h0;
  assign T_6150 = T_6148 | T_1782_26;
  assign T_6152 = T_1443 == 1'h0;
  assign T_6154 = T_6152 | T_1782_14;
  assign T_6156 = T_1380 == 1'h0;
  assign T_6158 = T_6156 | T_1782_7;
  assign T_6160 = T_1731 == 1'h0;
  assign T_6162 = T_6160 | T_1782_46;
  assign T_6164 = T_1596 == 1'h0;
  assign T_6166 = T_6164 | T_1782_31;
  assign T_6168 = T_1542 == 1'h0;
  assign T_6170 = T_6168 | T_1782_25;
  assign T_6172 = T_1695 == 1'h0;
  assign T_6174 = T_6172 | T_1782_42;
  assign T_6176 = T_1758 == 1'h0;
  assign T_6178 = T_6176 | T_1782_49;
  assign T_6442_0 = T_5880;
  assign T_6442_1 = 1'h1;
  assign T_6442_2 = T_5887;
  assign T_6442_3 = T_5891;
  assign T_6442_4 = T_5895;
  assign T_6442_5 = 1'h1;
  assign T_6442_6 = T_5902;
  assign T_6442_7 = T_5906;
  assign T_6442_8 = T_5910;
  assign T_6442_9 = 1'h1;
  assign T_6442_10 = 1'h1;
  assign T_6442_11 = 1'h1;
  assign T_6442_12 = 1'h1;
  assign T_6442_13 = 1'h1;
  assign T_6442_14 = 1'h1;
  assign T_6442_15 = 1'h1;
  assign T_6442_16 = T_5935;
  assign T_6442_17 = 1'h1;
  assign T_6442_18 = T_5942;
  assign T_6442_19 = T_5946;
  assign T_6442_20 = T_5950;
  assign T_6442_21 = 1'h1;
  assign T_6442_22 = T_5957;
  assign T_6442_23 = T_5961;
  assign T_6442_24 = T_5965;
  assign T_6442_25 = 1'h1;
  assign T_6442_26 = 1'h1;
  assign T_6442_27 = 1'h1;
  assign T_6442_28 = 1'h1;
  assign T_6442_29 = 1'h1;
  assign T_6442_30 = 1'h1;
  assign T_6442_31 = 1'h1;
  assign T_6442_32 = T_5990;
  assign T_6442_33 = T_5994;
  assign T_6442_34 = T_5998;
  assign T_6442_35 = T_6002;
  assign T_6442_36 = T_6006;
  assign T_6442_37 = T_6010;
  assign T_6442_38 = T_6014;
  assign T_6442_39 = T_6018;
  assign T_6442_40 = T_6022;
  assign T_6442_41 = T_6026;
  assign T_6442_42 = T_6030;
  assign T_6442_43 = T_6034;
  assign T_6442_44 = T_6038;
  assign T_6442_45 = T_6042;
  assign T_6442_46 = T_6046;
  assign T_6442_47 = T_6050;
  assign T_6442_48 = 1'h1;
  assign T_6442_49 = 1'h1;
  assign T_6442_50 = 1'h1;
  assign T_6442_51 = 1'h1;
  assign T_6442_52 = 1'h1;
  assign T_6442_53 = 1'h1;
  assign T_6442_54 = 1'h1;
  assign T_6442_55 = 1'h1;
  assign T_6442_56 = 1'h1;
  assign T_6442_57 = 1'h1;
  assign T_6442_58 = 1'h1;
  assign T_6442_59 = 1'h1;
  assign T_6442_60 = 1'h1;
  assign T_6442_61 = 1'h1;
  assign T_6442_62 = 1'h1;
  assign T_6442_63 = 1'h1;
  assign T_6442_64 = T_6102;
  assign T_6442_65 = T_6106;
  assign T_6442_66 = T_6110;
  assign T_6442_67 = T_6114;
  assign T_6442_68 = T_6118;
  assign T_6442_69 = T_6122;
  assign T_6442_70 = T_6126;
  assign T_6442_71 = T_6130;
  assign T_6442_72 = T_6134;
  assign T_6442_73 = T_6138;
  assign T_6442_74 = T_6142;
  assign T_6442_75 = T_6146;
  assign T_6442_76 = T_6150;
  assign T_6442_77 = T_6154;
  assign T_6442_78 = T_6158;
  assign T_6442_79 = T_6162;
  assign T_6442_80 = T_6166;
  assign T_6442_81 = T_6170;
  assign T_6442_82 = T_6174;
  assign T_6442_83 = T_6178;
  assign T_6442_84 = 1'h1;
  assign T_6442_85 = 1'h1;
  assign T_6442_86 = 1'h1;
  assign T_6442_87 = 1'h1;
  assign T_6442_88 = 1'h1;
  assign T_6442_89 = 1'h1;
  assign T_6442_90 = 1'h1;
  assign T_6442_91 = 1'h1;
  assign T_6442_92 = 1'h1;
  assign T_6442_93 = 1'h1;
  assign T_6442_94 = 1'h1;
  assign T_6442_95 = 1'h1;
  assign T_6442_96 = 1'h1;
  assign T_6442_97 = 1'h1;
  assign T_6442_98 = 1'h1;
  assign T_6442_99 = 1'h1;
  assign T_6442_100 = 1'h1;
  assign T_6442_101 = 1'h1;
  assign T_6442_102 = 1'h1;
  assign T_6442_103 = 1'h1;
  assign T_6442_104 = 1'h1;
  assign T_6442_105 = 1'h1;
  assign T_6442_106 = 1'h1;
  assign T_6442_107 = 1'h1;
  assign T_6442_108 = 1'h1;
  assign T_6442_109 = 1'h1;
  assign T_6442_110 = 1'h1;
  assign T_6442_111 = 1'h1;
  assign T_6442_112 = 1'h1;
  assign T_6442_113 = 1'h1;
  assign T_6442_114 = 1'h1;
  assign T_6442_115 = 1'h1;
  assign T_6442_116 = 1'h1;
  assign T_6442_117 = 1'h1;
  assign T_6442_118 = 1'h1;
  assign T_6442_119 = 1'h1;
  assign T_6442_120 = 1'h1;
  assign T_6442_121 = 1'h1;
  assign T_6442_122 = 1'h1;
  assign T_6442_123 = 1'h1;
  assign T_6442_124 = 1'h1;
  assign T_6442_125 = 1'h1;
  assign T_6442_126 = 1'h1;
  assign T_6442_127 = 1'h1;
  assign T_6576 = T_5878 | T_1787_1;
  assign T_6583 = T_5885 | T_1787_17;
  assign T_6587 = T_5889 | T_1787_30;
  assign T_6591 = T_5893 | T_1787_45;
  assign T_6598 = T_5900 | T_1787_9;
  assign T_6602 = T_5904 | T_1787_27;
  assign T_6606 = T_5908 | T_1787_40;
  assign T_6631 = T_5933 | T_1787_35;
  assign T_6638 = T_5940 | T_1787_33;
  assign T_6642 = T_5944 | T_1787_44;
  assign T_6646 = T_5948 | T_1787_5;
  assign T_6653 = T_5955 | T_1787_22;
  assign T_6657 = T_5959 | T_1787_39;
  assign T_6661 = T_5963 | T_1787_3;
  assign T_6686 = T_5988 | T_1787_18;
  assign T_6690 = T_5992 | T_1787_12;
  assign T_6694 = T_5996 | T_1787_19;
  assign T_6698 = T_6000 | T_1787_32;
  assign T_6702 = T_6004 | T_1787_43;
  assign T_6706 = T_6008 | T_1787_4;
  assign T_6710 = T_6012 | T_1787_10;
  assign T_6714 = T_6016 | T_1787_28;
  assign T_6718 = T_6020 | T_1787_38;
  assign T_6722 = T_6024 | T_1787_15;
  assign T_6726 = T_6028 | T_1787_2;
  assign T_6730 = T_6032 | T_1787_37;
  assign T_6734 = T_6036 | T_1787_23;
  assign T_6738 = T_6040 | T_1787_20;
  assign T_6742 = T_6044 | T_1787_6;
  assign T_6746 = T_6048 | T_1787_47;
  assign T_6798 = T_6100 | T_1787_21;
  assign T_6802 = T_6104 | T_1787_13;
  assign T_6806 = T_6108 | T_1787_29;
  assign T_6810 = T_6112 | T_1787_34;
  assign T_6814 = T_6116 | T_1787_48;
  assign T_6818 = T_6120 | T_1787_0;
  assign T_6822 = T_6124 | T_1787_11;
  assign T_6826 = T_6128 | T_1787_24;
  assign T_6830 = T_6132 | T_1787_36;
  assign T_6834 = T_6136 | T_1787_16;
  assign T_6838 = T_6140 | T_1787_8;
  assign T_6842 = T_6144 | T_1787_41;
  assign T_6846 = T_6148 | T_1787_26;
  assign T_6850 = T_6152 | T_1787_14;
  assign T_6854 = T_6156 | T_1787_7;
  assign T_6858 = T_6160 | T_1787_46;
  assign T_6862 = T_6164 | T_1787_31;
  assign T_6866 = T_6168 | T_1787_25;
  assign T_6870 = T_6172 | T_1787_42;
  assign T_6874 = T_6176 | T_1787_49;
  assign T_7138_0 = T_6576;
  assign T_7138_1 = 1'h1;
  assign T_7138_2 = T_6583;
  assign T_7138_3 = T_6587;
  assign T_7138_4 = T_6591;
  assign T_7138_5 = 1'h1;
  assign T_7138_6 = T_6598;
  assign T_7138_7 = T_6602;
  assign T_7138_8 = T_6606;
  assign T_7138_9 = 1'h1;
  assign T_7138_10 = 1'h1;
  assign T_7138_11 = 1'h1;
  assign T_7138_12 = 1'h1;
  assign T_7138_13 = 1'h1;
  assign T_7138_14 = 1'h1;
  assign T_7138_15 = 1'h1;
  assign T_7138_16 = T_6631;
  assign T_7138_17 = 1'h1;
  assign T_7138_18 = T_6638;
  assign T_7138_19 = T_6642;
  assign T_7138_20 = T_6646;
  assign T_7138_21 = 1'h1;
  assign T_7138_22 = T_6653;
  assign T_7138_23 = T_6657;
  assign T_7138_24 = T_6661;
  assign T_7138_25 = 1'h1;
  assign T_7138_26 = 1'h1;
  assign T_7138_27 = 1'h1;
  assign T_7138_28 = 1'h1;
  assign T_7138_29 = 1'h1;
  assign T_7138_30 = 1'h1;
  assign T_7138_31 = 1'h1;
  assign T_7138_32 = T_6686;
  assign T_7138_33 = T_6690;
  assign T_7138_34 = T_6694;
  assign T_7138_35 = T_6698;
  assign T_7138_36 = T_6702;
  assign T_7138_37 = T_6706;
  assign T_7138_38 = T_6710;
  assign T_7138_39 = T_6714;
  assign T_7138_40 = T_6718;
  assign T_7138_41 = T_6722;
  assign T_7138_42 = T_6726;
  assign T_7138_43 = T_6730;
  assign T_7138_44 = T_6734;
  assign T_7138_45 = T_6738;
  assign T_7138_46 = T_6742;
  assign T_7138_47 = T_6746;
  assign T_7138_48 = 1'h1;
  assign T_7138_49 = 1'h1;
  assign T_7138_50 = 1'h1;
  assign T_7138_51 = 1'h1;
  assign T_7138_52 = 1'h1;
  assign T_7138_53 = 1'h1;
  assign T_7138_54 = 1'h1;
  assign T_7138_55 = 1'h1;
  assign T_7138_56 = 1'h1;
  assign T_7138_57 = 1'h1;
  assign T_7138_58 = 1'h1;
  assign T_7138_59 = 1'h1;
  assign T_7138_60 = 1'h1;
  assign T_7138_61 = 1'h1;
  assign T_7138_62 = 1'h1;
  assign T_7138_63 = 1'h1;
  assign T_7138_64 = T_6798;
  assign T_7138_65 = T_6802;
  assign T_7138_66 = T_6806;
  assign T_7138_67 = T_6810;
  assign T_7138_68 = T_6814;
  assign T_7138_69 = T_6818;
  assign T_7138_70 = T_6822;
  assign T_7138_71 = T_6826;
  assign T_7138_72 = T_6830;
  assign T_7138_73 = T_6834;
  assign T_7138_74 = T_6838;
  assign T_7138_75 = T_6842;
  assign T_7138_76 = T_6846;
  assign T_7138_77 = T_6850;
  assign T_7138_78 = T_6854;
  assign T_7138_79 = T_6858;
  assign T_7138_80 = T_6862;
  assign T_7138_81 = T_6866;
  assign T_7138_82 = T_6870;
  assign T_7138_83 = T_6874;
  assign T_7138_84 = 1'h1;
  assign T_7138_85 = 1'h1;
  assign T_7138_86 = 1'h1;
  assign T_7138_87 = 1'h1;
  assign T_7138_88 = 1'h1;
  assign T_7138_89 = 1'h1;
  assign T_7138_90 = 1'h1;
  assign T_7138_91 = 1'h1;
  assign T_7138_92 = 1'h1;
  assign T_7138_93 = 1'h1;
  assign T_7138_94 = 1'h1;
  assign T_7138_95 = 1'h1;
  assign T_7138_96 = 1'h1;
  assign T_7138_97 = 1'h1;
  assign T_7138_98 = 1'h1;
  assign T_7138_99 = 1'h1;
  assign T_7138_100 = 1'h1;
  assign T_7138_101 = 1'h1;
  assign T_7138_102 = 1'h1;
  assign T_7138_103 = 1'h1;
  assign T_7138_104 = 1'h1;
  assign T_7138_105 = 1'h1;
  assign T_7138_106 = 1'h1;
  assign T_7138_107 = 1'h1;
  assign T_7138_108 = 1'h1;
  assign T_7138_109 = 1'h1;
  assign T_7138_110 = 1'h1;
  assign T_7138_111 = 1'h1;
  assign T_7138_112 = 1'h1;
  assign T_7138_113 = 1'h1;
  assign T_7138_114 = 1'h1;
  assign T_7138_115 = 1'h1;
  assign T_7138_116 = 1'h1;
  assign T_7138_117 = 1'h1;
  assign T_7138_118 = 1'h1;
  assign T_7138_119 = 1'h1;
  assign T_7138_120 = 1'h1;
  assign T_7138_121 = 1'h1;
  assign T_7138_122 = 1'h1;
  assign T_7138_123 = 1'h1;
  assign T_7138_124 = 1'h1;
  assign T_7138_125 = 1'h1;
  assign T_7138_126 = 1'h1;
  assign T_7138_127 = 1'h1;
  assign T_7269 = T_1028_bits_index[0];
  assign T_7270 = T_1028_bits_index[1];
  assign T_7271 = T_1028_bits_index[2];
  assign T_7272 = T_1028_bits_index[3];
  assign T_7273 = T_1028_bits_index[4];
  assign T_7274 = T_1028_bits_index[5];
  assign T_7275 = T_1028_bits_index[6];
  assign T_7279 = {T_7271,T_7270};
  assign T_7280 = {T_7279,T_7269};
  assign T_7281 = {T_7273,T_7272};
  assign T_7282 = {T_7275,T_7274};
  assign T_7283 = {T_7282,T_7281};
  assign T_7284 = {T_7283,T_7280};
  assign T_7285 = Queue_1_io_deq_bits_index[0];
  assign T_7286 = Queue_1_io_deq_bits_index[1];
  assign T_7287 = Queue_1_io_deq_bits_index[2];
  assign T_7288 = Queue_1_io_deq_bits_index[3];
  assign T_7289 = Queue_1_io_deq_bits_index[4];
  assign T_7290 = Queue_1_io_deq_bits_index[5];
  assign T_7291 = Queue_1_io_deq_bits_index[6];
  assign T_7295 = {T_7287,T_7286};
  assign T_7296 = {T_7295,T_7285};
  assign T_7297 = {T_7289,T_7288};
  assign T_7298 = {T_7291,T_7290};
  assign T_7299 = {T_7298,T_7297};
  assign T_7300 = {T_7299,T_7296};
  assign GEN_0 = GEN_148;
  assign GEN_22 = 7'h1 == T_7284 ? T_5050_1 : T_5050_0;
  assign GEN_23 = 7'h2 == T_7284 ? T_5050_2 : GEN_22;
  assign GEN_24 = 7'h3 == T_7284 ? T_5050_3 : GEN_23;
  assign GEN_25 = 7'h4 == T_7284 ? T_5050_4 : GEN_24;
  assign GEN_26 = 7'h5 == T_7284 ? T_5050_5 : GEN_25;
  assign GEN_27 = 7'h6 == T_7284 ? T_5050_6 : GEN_26;
  assign GEN_28 = 7'h7 == T_7284 ? T_5050_7 : GEN_27;
  assign GEN_29 = 7'h8 == T_7284 ? T_5050_8 : GEN_28;
  assign GEN_30 = 7'h9 == T_7284 ? T_5050_9 : GEN_29;
  assign GEN_31 = 7'ha == T_7284 ? T_5050_10 : GEN_30;
  assign GEN_32 = 7'hb == T_7284 ? T_5050_11 : GEN_31;
  assign GEN_33 = 7'hc == T_7284 ? T_5050_12 : GEN_32;
  assign GEN_34 = 7'hd == T_7284 ? T_5050_13 : GEN_33;
  assign GEN_35 = 7'he == T_7284 ? T_5050_14 : GEN_34;
  assign GEN_36 = 7'hf == T_7284 ? T_5050_15 : GEN_35;
  assign GEN_37 = 7'h10 == T_7284 ? T_5050_16 : GEN_36;
  assign GEN_38 = 7'h11 == T_7284 ? T_5050_17 : GEN_37;
  assign GEN_39 = 7'h12 == T_7284 ? T_5050_18 : GEN_38;
  assign GEN_40 = 7'h13 == T_7284 ? T_5050_19 : GEN_39;
  assign GEN_41 = 7'h14 == T_7284 ? T_5050_20 : GEN_40;
  assign GEN_42 = 7'h15 == T_7284 ? T_5050_21 : GEN_41;
  assign GEN_43 = 7'h16 == T_7284 ? T_5050_22 : GEN_42;
  assign GEN_44 = 7'h17 == T_7284 ? T_5050_23 : GEN_43;
  assign GEN_45 = 7'h18 == T_7284 ? T_5050_24 : GEN_44;
  assign GEN_46 = 7'h19 == T_7284 ? T_5050_25 : GEN_45;
  assign GEN_47 = 7'h1a == T_7284 ? T_5050_26 : GEN_46;
  assign GEN_48 = 7'h1b == T_7284 ? T_5050_27 : GEN_47;
  assign GEN_49 = 7'h1c == T_7284 ? T_5050_28 : GEN_48;
  assign GEN_50 = 7'h1d == T_7284 ? T_5050_29 : GEN_49;
  assign GEN_51 = 7'h1e == T_7284 ? T_5050_30 : GEN_50;
  assign GEN_52 = 7'h1f == T_7284 ? T_5050_31 : GEN_51;
  assign GEN_53 = 7'h20 == T_7284 ? T_5050_32 : GEN_52;
  assign GEN_54 = 7'h21 == T_7284 ? T_5050_33 : GEN_53;
  assign GEN_55 = 7'h22 == T_7284 ? T_5050_34 : GEN_54;
  assign GEN_56 = 7'h23 == T_7284 ? T_5050_35 : GEN_55;
  assign GEN_57 = 7'h24 == T_7284 ? T_5050_36 : GEN_56;
  assign GEN_58 = 7'h25 == T_7284 ? T_5050_37 : GEN_57;
  assign GEN_59 = 7'h26 == T_7284 ? T_5050_38 : GEN_58;
  assign GEN_60 = 7'h27 == T_7284 ? T_5050_39 : GEN_59;
  assign GEN_61 = 7'h28 == T_7284 ? T_5050_40 : GEN_60;
  assign GEN_62 = 7'h29 == T_7284 ? T_5050_41 : GEN_61;
  assign GEN_63 = 7'h2a == T_7284 ? T_5050_42 : GEN_62;
  assign GEN_64 = 7'h2b == T_7284 ? T_5050_43 : GEN_63;
  assign GEN_65 = 7'h2c == T_7284 ? T_5050_44 : GEN_64;
  assign GEN_66 = 7'h2d == T_7284 ? T_5050_45 : GEN_65;
  assign GEN_67 = 7'h2e == T_7284 ? T_5050_46 : GEN_66;
  assign GEN_68 = 7'h2f == T_7284 ? T_5050_47 : GEN_67;
  assign GEN_69 = 7'h30 == T_7284 ? T_5050_48 : GEN_68;
  assign GEN_70 = 7'h31 == T_7284 ? T_5050_49 : GEN_69;
  assign GEN_71 = 7'h32 == T_7284 ? T_5050_50 : GEN_70;
  assign GEN_72 = 7'h33 == T_7284 ? T_5050_51 : GEN_71;
  assign GEN_73 = 7'h34 == T_7284 ? T_5050_52 : GEN_72;
  assign GEN_74 = 7'h35 == T_7284 ? T_5050_53 : GEN_73;
  assign GEN_75 = 7'h36 == T_7284 ? T_5050_54 : GEN_74;
  assign GEN_76 = 7'h37 == T_7284 ? T_5050_55 : GEN_75;
  assign GEN_77 = 7'h38 == T_7284 ? T_5050_56 : GEN_76;
  assign GEN_78 = 7'h39 == T_7284 ? T_5050_57 : GEN_77;
  assign GEN_79 = 7'h3a == T_7284 ? T_5050_58 : GEN_78;
  assign GEN_80 = 7'h3b == T_7284 ? T_5050_59 : GEN_79;
  assign GEN_81 = 7'h3c == T_7284 ? T_5050_60 : GEN_80;
  assign GEN_82 = 7'h3d == T_7284 ? T_5050_61 : GEN_81;
  assign GEN_83 = 7'h3e == T_7284 ? T_5050_62 : GEN_82;
  assign GEN_84 = 7'h3f == T_7284 ? T_5050_63 : GEN_83;
  assign GEN_85 = 7'h40 == T_7284 ? T_5050_64 : GEN_84;
  assign GEN_86 = 7'h41 == T_7284 ? T_5050_65 : GEN_85;
  assign GEN_87 = 7'h42 == T_7284 ? T_5050_66 : GEN_86;
  assign GEN_88 = 7'h43 == T_7284 ? T_5050_67 : GEN_87;
  assign GEN_89 = 7'h44 == T_7284 ? T_5050_68 : GEN_88;
  assign GEN_90 = 7'h45 == T_7284 ? T_5050_69 : GEN_89;
  assign GEN_91 = 7'h46 == T_7284 ? T_5050_70 : GEN_90;
  assign GEN_92 = 7'h47 == T_7284 ? T_5050_71 : GEN_91;
  assign GEN_93 = 7'h48 == T_7284 ? T_5050_72 : GEN_92;
  assign GEN_94 = 7'h49 == T_7284 ? T_5050_73 : GEN_93;
  assign GEN_95 = 7'h4a == T_7284 ? T_5050_74 : GEN_94;
  assign GEN_96 = 7'h4b == T_7284 ? T_5050_75 : GEN_95;
  assign GEN_97 = 7'h4c == T_7284 ? T_5050_76 : GEN_96;
  assign GEN_98 = 7'h4d == T_7284 ? T_5050_77 : GEN_97;
  assign GEN_99 = 7'h4e == T_7284 ? T_5050_78 : GEN_98;
  assign GEN_100 = 7'h4f == T_7284 ? T_5050_79 : GEN_99;
  assign GEN_101 = 7'h50 == T_7284 ? T_5050_80 : GEN_100;
  assign GEN_102 = 7'h51 == T_7284 ? T_5050_81 : GEN_101;
  assign GEN_103 = 7'h52 == T_7284 ? T_5050_82 : GEN_102;
  assign GEN_104 = 7'h53 == T_7284 ? T_5050_83 : GEN_103;
  assign GEN_105 = 7'h54 == T_7284 ? T_5050_84 : GEN_104;
  assign GEN_106 = 7'h55 == T_7284 ? T_5050_85 : GEN_105;
  assign GEN_107 = 7'h56 == T_7284 ? T_5050_86 : GEN_106;
  assign GEN_108 = 7'h57 == T_7284 ? T_5050_87 : GEN_107;
  assign GEN_109 = 7'h58 == T_7284 ? T_5050_88 : GEN_108;
  assign GEN_110 = 7'h59 == T_7284 ? T_5050_89 : GEN_109;
  assign GEN_111 = 7'h5a == T_7284 ? T_5050_90 : GEN_110;
  assign GEN_112 = 7'h5b == T_7284 ? T_5050_91 : GEN_111;
  assign GEN_113 = 7'h5c == T_7284 ? T_5050_92 : GEN_112;
  assign GEN_114 = 7'h5d == T_7284 ? T_5050_93 : GEN_113;
  assign GEN_115 = 7'h5e == T_7284 ? T_5050_94 : GEN_114;
  assign GEN_116 = 7'h5f == T_7284 ? T_5050_95 : GEN_115;
  assign GEN_117 = 7'h60 == T_7284 ? T_5050_96 : GEN_116;
  assign GEN_118 = 7'h61 == T_7284 ? T_5050_97 : GEN_117;
  assign GEN_119 = 7'h62 == T_7284 ? T_5050_98 : GEN_118;
  assign GEN_120 = 7'h63 == T_7284 ? T_5050_99 : GEN_119;
  assign GEN_121 = 7'h64 == T_7284 ? T_5050_100 : GEN_120;
  assign GEN_122 = 7'h65 == T_7284 ? T_5050_101 : GEN_121;
  assign GEN_123 = 7'h66 == T_7284 ? T_5050_102 : GEN_122;
  assign GEN_124 = 7'h67 == T_7284 ? T_5050_103 : GEN_123;
  assign GEN_125 = 7'h68 == T_7284 ? T_5050_104 : GEN_124;
  assign GEN_126 = 7'h69 == T_7284 ? T_5050_105 : GEN_125;
  assign GEN_127 = 7'h6a == T_7284 ? T_5050_106 : GEN_126;
  assign GEN_128 = 7'h6b == T_7284 ? T_5050_107 : GEN_127;
  assign GEN_129 = 7'h6c == T_7284 ? T_5050_108 : GEN_128;
  assign GEN_130 = 7'h6d == T_7284 ? T_5050_109 : GEN_129;
  assign GEN_131 = 7'h6e == T_7284 ? T_5050_110 : GEN_130;
  assign GEN_132 = 7'h6f == T_7284 ? T_5050_111 : GEN_131;
  assign GEN_133 = 7'h70 == T_7284 ? T_5050_112 : GEN_132;
  assign GEN_134 = 7'h71 == T_7284 ? T_5050_113 : GEN_133;
  assign GEN_135 = 7'h72 == T_7284 ? T_5050_114 : GEN_134;
  assign GEN_136 = 7'h73 == T_7284 ? T_5050_115 : GEN_135;
  assign GEN_137 = 7'h74 == T_7284 ? T_5050_116 : GEN_136;
  assign GEN_138 = 7'h75 == T_7284 ? T_5050_117 : GEN_137;
  assign GEN_139 = 7'h76 == T_7284 ? T_5050_118 : GEN_138;
  assign GEN_140 = 7'h77 == T_7284 ? T_5050_119 : GEN_139;
  assign GEN_141 = 7'h78 == T_7284 ? T_5050_120 : GEN_140;
  assign GEN_142 = 7'h79 == T_7284 ? T_5050_121 : GEN_141;
  assign GEN_143 = 7'h7a == T_7284 ? T_5050_122 : GEN_142;
  assign GEN_144 = 7'h7b == T_7284 ? T_5050_123 : GEN_143;
  assign GEN_145 = 7'h7c == T_7284 ? T_5050_124 : GEN_144;
  assign GEN_146 = 7'h7d == T_7284 ? T_5050_125 : GEN_145;
  assign GEN_147 = 7'h7e == T_7284 ? T_5050_126 : GEN_146;
  assign GEN_148 = 7'h7f == T_7284 ? T_5050_127 : GEN_147;
  assign GEN_1 = GEN_275;
  assign GEN_149 = 7'h1 == T_7284 ? T_5746_1 : T_5746_0;
  assign GEN_150 = 7'h2 == T_7284 ? T_5746_2 : GEN_149;
  assign GEN_151 = 7'h3 == T_7284 ? T_5746_3 : GEN_150;
  assign GEN_152 = 7'h4 == T_7284 ? T_5746_4 : GEN_151;
  assign GEN_153 = 7'h5 == T_7284 ? T_5746_5 : GEN_152;
  assign GEN_154 = 7'h6 == T_7284 ? T_5746_6 : GEN_153;
  assign GEN_155 = 7'h7 == T_7284 ? T_5746_7 : GEN_154;
  assign GEN_156 = 7'h8 == T_7284 ? T_5746_8 : GEN_155;
  assign GEN_157 = 7'h9 == T_7284 ? T_5746_9 : GEN_156;
  assign GEN_158 = 7'ha == T_7284 ? T_5746_10 : GEN_157;
  assign GEN_159 = 7'hb == T_7284 ? T_5746_11 : GEN_158;
  assign GEN_160 = 7'hc == T_7284 ? T_5746_12 : GEN_159;
  assign GEN_161 = 7'hd == T_7284 ? T_5746_13 : GEN_160;
  assign GEN_162 = 7'he == T_7284 ? T_5746_14 : GEN_161;
  assign GEN_163 = 7'hf == T_7284 ? T_5746_15 : GEN_162;
  assign GEN_164 = 7'h10 == T_7284 ? T_5746_16 : GEN_163;
  assign GEN_165 = 7'h11 == T_7284 ? T_5746_17 : GEN_164;
  assign GEN_166 = 7'h12 == T_7284 ? T_5746_18 : GEN_165;
  assign GEN_167 = 7'h13 == T_7284 ? T_5746_19 : GEN_166;
  assign GEN_168 = 7'h14 == T_7284 ? T_5746_20 : GEN_167;
  assign GEN_169 = 7'h15 == T_7284 ? T_5746_21 : GEN_168;
  assign GEN_170 = 7'h16 == T_7284 ? T_5746_22 : GEN_169;
  assign GEN_171 = 7'h17 == T_7284 ? T_5746_23 : GEN_170;
  assign GEN_172 = 7'h18 == T_7284 ? T_5746_24 : GEN_171;
  assign GEN_173 = 7'h19 == T_7284 ? T_5746_25 : GEN_172;
  assign GEN_174 = 7'h1a == T_7284 ? T_5746_26 : GEN_173;
  assign GEN_175 = 7'h1b == T_7284 ? T_5746_27 : GEN_174;
  assign GEN_176 = 7'h1c == T_7284 ? T_5746_28 : GEN_175;
  assign GEN_177 = 7'h1d == T_7284 ? T_5746_29 : GEN_176;
  assign GEN_178 = 7'h1e == T_7284 ? T_5746_30 : GEN_177;
  assign GEN_179 = 7'h1f == T_7284 ? T_5746_31 : GEN_178;
  assign GEN_180 = 7'h20 == T_7284 ? T_5746_32 : GEN_179;
  assign GEN_181 = 7'h21 == T_7284 ? T_5746_33 : GEN_180;
  assign GEN_182 = 7'h22 == T_7284 ? T_5746_34 : GEN_181;
  assign GEN_183 = 7'h23 == T_7284 ? T_5746_35 : GEN_182;
  assign GEN_184 = 7'h24 == T_7284 ? T_5746_36 : GEN_183;
  assign GEN_185 = 7'h25 == T_7284 ? T_5746_37 : GEN_184;
  assign GEN_186 = 7'h26 == T_7284 ? T_5746_38 : GEN_185;
  assign GEN_187 = 7'h27 == T_7284 ? T_5746_39 : GEN_186;
  assign GEN_188 = 7'h28 == T_7284 ? T_5746_40 : GEN_187;
  assign GEN_189 = 7'h29 == T_7284 ? T_5746_41 : GEN_188;
  assign GEN_190 = 7'h2a == T_7284 ? T_5746_42 : GEN_189;
  assign GEN_191 = 7'h2b == T_7284 ? T_5746_43 : GEN_190;
  assign GEN_192 = 7'h2c == T_7284 ? T_5746_44 : GEN_191;
  assign GEN_193 = 7'h2d == T_7284 ? T_5746_45 : GEN_192;
  assign GEN_194 = 7'h2e == T_7284 ? T_5746_46 : GEN_193;
  assign GEN_195 = 7'h2f == T_7284 ? T_5746_47 : GEN_194;
  assign GEN_196 = 7'h30 == T_7284 ? T_5746_48 : GEN_195;
  assign GEN_197 = 7'h31 == T_7284 ? T_5746_49 : GEN_196;
  assign GEN_198 = 7'h32 == T_7284 ? T_5746_50 : GEN_197;
  assign GEN_199 = 7'h33 == T_7284 ? T_5746_51 : GEN_198;
  assign GEN_200 = 7'h34 == T_7284 ? T_5746_52 : GEN_199;
  assign GEN_201 = 7'h35 == T_7284 ? T_5746_53 : GEN_200;
  assign GEN_202 = 7'h36 == T_7284 ? T_5746_54 : GEN_201;
  assign GEN_203 = 7'h37 == T_7284 ? T_5746_55 : GEN_202;
  assign GEN_204 = 7'h38 == T_7284 ? T_5746_56 : GEN_203;
  assign GEN_205 = 7'h39 == T_7284 ? T_5746_57 : GEN_204;
  assign GEN_206 = 7'h3a == T_7284 ? T_5746_58 : GEN_205;
  assign GEN_207 = 7'h3b == T_7284 ? T_5746_59 : GEN_206;
  assign GEN_208 = 7'h3c == T_7284 ? T_5746_60 : GEN_207;
  assign GEN_209 = 7'h3d == T_7284 ? T_5746_61 : GEN_208;
  assign GEN_210 = 7'h3e == T_7284 ? T_5746_62 : GEN_209;
  assign GEN_211 = 7'h3f == T_7284 ? T_5746_63 : GEN_210;
  assign GEN_212 = 7'h40 == T_7284 ? T_5746_64 : GEN_211;
  assign GEN_213 = 7'h41 == T_7284 ? T_5746_65 : GEN_212;
  assign GEN_214 = 7'h42 == T_7284 ? T_5746_66 : GEN_213;
  assign GEN_215 = 7'h43 == T_7284 ? T_5746_67 : GEN_214;
  assign GEN_216 = 7'h44 == T_7284 ? T_5746_68 : GEN_215;
  assign GEN_217 = 7'h45 == T_7284 ? T_5746_69 : GEN_216;
  assign GEN_218 = 7'h46 == T_7284 ? T_5746_70 : GEN_217;
  assign GEN_219 = 7'h47 == T_7284 ? T_5746_71 : GEN_218;
  assign GEN_220 = 7'h48 == T_7284 ? T_5746_72 : GEN_219;
  assign GEN_221 = 7'h49 == T_7284 ? T_5746_73 : GEN_220;
  assign GEN_222 = 7'h4a == T_7284 ? T_5746_74 : GEN_221;
  assign GEN_223 = 7'h4b == T_7284 ? T_5746_75 : GEN_222;
  assign GEN_224 = 7'h4c == T_7284 ? T_5746_76 : GEN_223;
  assign GEN_225 = 7'h4d == T_7284 ? T_5746_77 : GEN_224;
  assign GEN_226 = 7'h4e == T_7284 ? T_5746_78 : GEN_225;
  assign GEN_227 = 7'h4f == T_7284 ? T_5746_79 : GEN_226;
  assign GEN_228 = 7'h50 == T_7284 ? T_5746_80 : GEN_227;
  assign GEN_229 = 7'h51 == T_7284 ? T_5746_81 : GEN_228;
  assign GEN_230 = 7'h52 == T_7284 ? T_5746_82 : GEN_229;
  assign GEN_231 = 7'h53 == T_7284 ? T_5746_83 : GEN_230;
  assign GEN_232 = 7'h54 == T_7284 ? T_5746_84 : GEN_231;
  assign GEN_233 = 7'h55 == T_7284 ? T_5746_85 : GEN_232;
  assign GEN_234 = 7'h56 == T_7284 ? T_5746_86 : GEN_233;
  assign GEN_235 = 7'h57 == T_7284 ? T_5746_87 : GEN_234;
  assign GEN_236 = 7'h58 == T_7284 ? T_5746_88 : GEN_235;
  assign GEN_237 = 7'h59 == T_7284 ? T_5746_89 : GEN_236;
  assign GEN_238 = 7'h5a == T_7284 ? T_5746_90 : GEN_237;
  assign GEN_239 = 7'h5b == T_7284 ? T_5746_91 : GEN_238;
  assign GEN_240 = 7'h5c == T_7284 ? T_5746_92 : GEN_239;
  assign GEN_241 = 7'h5d == T_7284 ? T_5746_93 : GEN_240;
  assign GEN_242 = 7'h5e == T_7284 ? T_5746_94 : GEN_241;
  assign GEN_243 = 7'h5f == T_7284 ? T_5746_95 : GEN_242;
  assign GEN_244 = 7'h60 == T_7284 ? T_5746_96 : GEN_243;
  assign GEN_245 = 7'h61 == T_7284 ? T_5746_97 : GEN_244;
  assign GEN_246 = 7'h62 == T_7284 ? T_5746_98 : GEN_245;
  assign GEN_247 = 7'h63 == T_7284 ? T_5746_99 : GEN_246;
  assign GEN_248 = 7'h64 == T_7284 ? T_5746_100 : GEN_247;
  assign GEN_249 = 7'h65 == T_7284 ? T_5746_101 : GEN_248;
  assign GEN_250 = 7'h66 == T_7284 ? T_5746_102 : GEN_249;
  assign GEN_251 = 7'h67 == T_7284 ? T_5746_103 : GEN_250;
  assign GEN_252 = 7'h68 == T_7284 ? T_5746_104 : GEN_251;
  assign GEN_253 = 7'h69 == T_7284 ? T_5746_105 : GEN_252;
  assign GEN_254 = 7'h6a == T_7284 ? T_5746_106 : GEN_253;
  assign GEN_255 = 7'h6b == T_7284 ? T_5746_107 : GEN_254;
  assign GEN_256 = 7'h6c == T_7284 ? T_5746_108 : GEN_255;
  assign GEN_257 = 7'h6d == T_7284 ? T_5746_109 : GEN_256;
  assign GEN_258 = 7'h6e == T_7284 ? T_5746_110 : GEN_257;
  assign GEN_259 = 7'h6f == T_7284 ? T_5746_111 : GEN_258;
  assign GEN_260 = 7'h70 == T_7284 ? T_5746_112 : GEN_259;
  assign GEN_261 = 7'h71 == T_7284 ? T_5746_113 : GEN_260;
  assign GEN_262 = 7'h72 == T_7284 ? T_5746_114 : GEN_261;
  assign GEN_263 = 7'h73 == T_7284 ? T_5746_115 : GEN_262;
  assign GEN_264 = 7'h74 == T_7284 ? T_5746_116 : GEN_263;
  assign GEN_265 = 7'h75 == T_7284 ? T_5746_117 : GEN_264;
  assign GEN_266 = 7'h76 == T_7284 ? T_5746_118 : GEN_265;
  assign GEN_267 = 7'h77 == T_7284 ? T_5746_119 : GEN_266;
  assign GEN_268 = 7'h78 == T_7284 ? T_5746_120 : GEN_267;
  assign GEN_269 = 7'h79 == T_7284 ? T_5746_121 : GEN_268;
  assign GEN_270 = 7'h7a == T_7284 ? T_5746_122 : GEN_269;
  assign GEN_271 = 7'h7b == T_7284 ? T_5746_123 : GEN_270;
  assign GEN_272 = 7'h7c == T_7284 ? T_5746_124 : GEN_271;
  assign GEN_273 = 7'h7d == T_7284 ? T_5746_125 : GEN_272;
  assign GEN_274 = 7'h7e == T_7284 ? T_5746_126 : GEN_273;
  assign GEN_275 = 7'h7f == T_7284 ? T_5746_127 : GEN_274;
  assign T_7303 = T_1028_bits_read ? GEN_0 : GEN_1;
  assign GEN_2 = GEN_402;
  assign GEN_276 = 7'h1 == T_7300 ? T_6442_1 : T_6442_0;
  assign GEN_277 = 7'h2 == T_7300 ? T_6442_2 : GEN_276;
  assign GEN_278 = 7'h3 == T_7300 ? T_6442_3 : GEN_277;
  assign GEN_279 = 7'h4 == T_7300 ? T_6442_4 : GEN_278;
  assign GEN_280 = 7'h5 == T_7300 ? T_6442_5 : GEN_279;
  assign GEN_281 = 7'h6 == T_7300 ? T_6442_6 : GEN_280;
  assign GEN_282 = 7'h7 == T_7300 ? T_6442_7 : GEN_281;
  assign GEN_283 = 7'h8 == T_7300 ? T_6442_8 : GEN_282;
  assign GEN_284 = 7'h9 == T_7300 ? T_6442_9 : GEN_283;
  assign GEN_285 = 7'ha == T_7300 ? T_6442_10 : GEN_284;
  assign GEN_286 = 7'hb == T_7300 ? T_6442_11 : GEN_285;
  assign GEN_287 = 7'hc == T_7300 ? T_6442_12 : GEN_286;
  assign GEN_288 = 7'hd == T_7300 ? T_6442_13 : GEN_287;
  assign GEN_289 = 7'he == T_7300 ? T_6442_14 : GEN_288;
  assign GEN_290 = 7'hf == T_7300 ? T_6442_15 : GEN_289;
  assign GEN_291 = 7'h10 == T_7300 ? T_6442_16 : GEN_290;
  assign GEN_292 = 7'h11 == T_7300 ? T_6442_17 : GEN_291;
  assign GEN_293 = 7'h12 == T_7300 ? T_6442_18 : GEN_292;
  assign GEN_294 = 7'h13 == T_7300 ? T_6442_19 : GEN_293;
  assign GEN_295 = 7'h14 == T_7300 ? T_6442_20 : GEN_294;
  assign GEN_296 = 7'h15 == T_7300 ? T_6442_21 : GEN_295;
  assign GEN_297 = 7'h16 == T_7300 ? T_6442_22 : GEN_296;
  assign GEN_298 = 7'h17 == T_7300 ? T_6442_23 : GEN_297;
  assign GEN_299 = 7'h18 == T_7300 ? T_6442_24 : GEN_298;
  assign GEN_300 = 7'h19 == T_7300 ? T_6442_25 : GEN_299;
  assign GEN_301 = 7'h1a == T_7300 ? T_6442_26 : GEN_300;
  assign GEN_302 = 7'h1b == T_7300 ? T_6442_27 : GEN_301;
  assign GEN_303 = 7'h1c == T_7300 ? T_6442_28 : GEN_302;
  assign GEN_304 = 7'h1d == T_7300 ? T_6442_29 : GEN_303;
  assign GEN_305 = 7'h1e == T_7300 ? T_6442_30 : GEN_304;
  assign GEN_306 = 7'h1f == T_7300 ? T_6442_31 : GEN_305;
  assign GEN_307 = 7'h20 == T_7300 ? T_6442_32 : GEN_306;
  assign GEN_308 = 7'h21 == T_7300 ? T_6442_33 : GEN_307;
  assign GEN_309 = 7'h22 == T_7300 ? T_6442_34 : GEN_308;
  assign GEN_310 = 7'h23 == T_7300 ? T_6442_35 : GEN_309;
  assign GEN_311 = 7'h24 == T_7300 ? T_6442_36 : GEN_310;
  assign GEN_312 = 7'h25 == T_7300 ? T_6442_37 : GEN_311;
  assign GEN_313 = 7'h26 == T_7300 ? T_6442_38 : GEN_312;
  assign GEN_314 = 7'h27 == T_7300 ? T_6442_39 : GEN_313;
  assign GEN_315 = 7'h28 == T_7300 ? T_6442_40 : GEN_314;
  assign GEN_316 = 7'h29 == T_7300 ? T_6442_41 : GEN_315;
  assign GEN_317 = 7'h2a == T_7300 ? T_6442_42 : GEN_316;
  assign GEN_318 = 7'h2b == T_7300 ? T_6442_43 : GEN_317;
  assign GEN_319 = 7'h2c == T_7300 ? T_6442_44 : GEN_318;
  assign GEN_320 = 7'h2d == T_7300 ? T_6442_45 : GEN_319;
  assign GEN_321 = 7'h2e == T_7300 ? T_6442_46 : GEN_320;
  assign GEN_322 = 7'h2f == T_7300 ? T_6442_47 : GEN_321;
  assign GEN_323 = 7'h30 == T_7300 ? T_6442_48 : GEN_322;
  assign GEN_324 = 7'h31 == T_7300 ? T_6442_49 : GEN_323;
  assign GEN_325 = 7'h32 == T_7300 ? T_6442_50 : GEN_324;
  assign GEN_326 = 7'h33 == T_7300 ? T_6442_51 : GEN_325;
  assign GEN_327 = 7'h34 == T_7300 ? T_6442_52 : GEN_326;
  assign GEN_328 = 7'h35 == T_7300 ? T_6442_53 : GEN_327;
  assign GEN_329 = 7'h36 == T_7300 ? T_6442_54 : GEN_328;
  assign GEN_330 = 7'h37 == T_7300 ? T_6442_55 : GEN_329;
  assign GEN_331 = 7'h38 == T_7300 ? T_6442_56 : GEN_330;
  assign GEN_332 = 7'h39 == T_7300 ? T_6442_57 : GEN_331;
  assign GEN_333 = 7'h3a == T_7300 ? T_6442_58 : GEN_332;
  assign GEN_334 = 7'h3b == T_7300 ? T_6442_59 : GEN_333;
  assign GEN_335 = 7'h3c == T_7300 ? T_6442_60 : GEN_334;
  assign GEN_336 = 7'h3d == T_7300 ? T_6442_61 : GEN_335;
  assign GEN_337 = 7'h3e == T_7300 ? T_6442_62 : GEN_336;
  assign GEN_338 = 7'h3f == T_7300 ? T_6442_63 : GEN_337;
  assign GEN_339 = 7'h40 == T_7300 ? T_6442_64 : GEN_338;
  assign GEN_340 = 7'h41 == T_7300 ? T_6442_65 : GEN_339;
  assign GEN_341 = 7'h42 == T_7300 ? T_6442_66 : GEN_340;
  assign GEN_342 = 7'h43 == T_7300 ? T_6442_67 : GEN_341;
  assign GEN_343 = 7'h44 == T_7300 ? T_6442_68 : GEN_342;
  assign GEN_344 = 7'h45 == T_7300 ? T_6442_69 : GEN_343;
  assign GEN_345 = 7'h46 == T_7300 ? T_6442_70 : GEN_344;
  assign GEN_346 = 7'h47 == T_7300 ? T_6442_71 : GEN_345;
  assign GEN_347 = 7'h48 == T_7300 ? T_6442_72 : GEN_346;
  assign GEN_348 = 7'h49 == T_7300 ? T_6442_73 : GEN_347;
  assign GEN_349 = 7'h4a == T_7300 ? T_6442_74 : GEN_348;
  assign GEN_350 = 7'h4b == T_7300 ? T_6442_75 : GEN_349;
  assign GEN_351 = 7'h4c == T_7300 ? T_6442_76 : GEN_350;
  assign GEN_352 = 7'h4d == T_7300 ? T_6442_77 : GEN_351;
  assign GEN_353 = 7'h4e == T_7300 ? T_6442_78 : GEN_352;
  assign GEN_354 = 7'h4f == T_7300 ? T_6442_79 : GEN_353;
  assign GEN_355 = 7'h50 == T_7300 ? T_6442_80 : GEN_354;
  assign GEN_356 = 7'h51 == T_7300 ? T_6442_81 : GEN_355;
  assign GEN_357 = 7'h52 == T_7300 ? T_6442_82 : GEN_356;
  assign GEN_358 = 7'h53 == T_7300 ? T_6442_83 : GEN_357;
  assign GEN_359 = 7'h54 == T_7300 ? T_6442_84 : GEN_358;
  assign GEN_360 = 7'h55 == T_7300 ? T_6442_85 : GEN_359;
  assign GEN_361 = 7'h56 == T_7300 ? T_6442_86 : GEN_360;
  assign GEN_362 = 7'h57 == T_7300 ? T_6442_87 : GEN_361;
  assign GEN_363 = 7'h58 == T_7300 ? T_6442_88 : GEN_362;
  assign GEN_364 = 7'h59 == T_7300 ? T_6442_89 : GEN_363;
  assign GEN_365 = 7'h5a == T_7300 ? T_6442_90 : GEN_364;
  assign GEN_366 = 7'h5b == T_7300 ? T_6442_91 : GEN_365;
  assign GEN_367 = 7'h5c == T_7300 ? T_6442_92 : GEN_366;
  assign GEN_368 = 7'h5d == T_7300 ? T_6442_93 : GEN_367;
  assign GEN_369 = 7'h5e == T_7300 ? T_6442_94 : GEN_368;
  assign GEN_370 = 7'h5f == T_7300 ? T_6442_95 : GEN_369;
  assign GEN_371 = 7'h60 == T_7300 ? T_6442_96 : GEN_370;
  assign GEN_372 = 7'h61 == T_7300 ? T_6442_97 : GEN_371;
  assign GEN_373 = 7'h62 == T_7300 ? T_6442_98 : GEN_372;
  assign GEN_374 = 7'h63 == T_7300 ? T_6442_99 : GEN_373;
  assign GEN_375 = 7'h64 == T_7300 ? T_6442_100 : GEN_374;
  assign GEN_376 = 7'h65 == T_7300 ? T_6442_101 : GEN_375;
  assign GEN_377 = 7'h66 == T_7300 ? T_6442_102 : GEN_376;
  assign GEN_378 = 7'h67 == T_7300 ? T_6442_103 : GEN_377;
  assign GEN_379 = 7'h68 == T_7300 ? T_6442_104 : GEN_378;
  assign GEN_380 = 7'h69 == T_7300 ? T_6442_105 : GEN_379;
  assign GEN_381 = 7'h6a == T_7300 ? T_6442_106 : GEN_380;
  assign GEN_382 = 7'h6b == T_7300 ? T_6442_107 : GEN_381;
  assign GEN_383 = 7'h6c == T_7300 ? T_6442_108 : GEN_382;
  assign GEN_384 = 7'h6d == T_7300 ? T_6442_109 : GEN_383;
  assign GEN_385 = 7'h6e == T_7300 ? T_6442_110 : GEN_384;
  assign GEN_386 = 7'h6f == T_7300 ? T_6442_111 : GEN_385;
  assign GEN_387 = 7'h70 == T_7300 ? T_6442_112 : GEN_386;
  assign GEN_388 = 7'h71 == T_7300 ? T_6442_113 : GEN_387;
  assign GEN_389 = 7'h72 == T_7300 ? T_6442_114 : GEN_388;
  assign GEN_390 = 7'h73 == T_7300 ? T_6442_115 : GEN_389;
  assign GEN_391 = 7'h74 == T_7300 ? T_6442_116 : GEN_390;
  assign GEN_392 = 7'h75 == T_7300 ? T_6442_117 : GEN_391;
  assign GEN_393 = 7'h76 == T_7300 ? T_6442_118 : GEN_392;
  assign GEN_394 = 7'h77 == T_7300 ? T_6442_119 : GEN_393;
  assign GEN_395 = 7'h78 == T_7300 ? T_6442_120 : GEN_394;
  assign GEN_396 = 7'h79 == T_7300 ? T_6442_121 : GEN_395;
  assign GEN_397 = 7'h7a == T_7300 ? T_6442_122 : GEN_396;
  assign GEN_398 = 7'h7b == T_7300 ? T_6442_123 : GEN_397;
  assign GEN_399 = 7'h7c == T_7300 ? T_6442_124 : GEN_398;
  assign GEN_400 = 7'h7d == T_7300 ? T_6442_125 : GEN_399;
  assign GEN_401 = 7'h7e == T_7300 ? T_6442_126 : GEN_400;
  assign GEN_402 = 7'h7f == T_7300 ? T_6442_127 : GEN_401;
  assign GEN_3 = GEN_529;
  assign GEN_403 = 7'h1 == T_7300 ? T_7138_1 : T_7138_0;
  assign GEN_404 = 7'h2 == T_7300 ? T_7138_2 : GEN_403;
  assign GEN_405 = 7'h3 == T_7300 ? T_7138_3 : GEN_404;
  assign GEN_406 = 7'h4 == T_7300 ? T_7138_4 : GEN_405;
  assign GEN_407 = 7'h5 == T_7300 ? T_7138_5 : GEN_406;
  assign GEN_408 = 7'h6 == T_7300 ? T_7138_6 : GEN_407;
  assign GEN_409 = 7'h7 == T_7300 ? T_7138_7 : GEN_408;
  assign GEN_410 = 7'h8 == T_7300 ? T_7138_8 : GEN_409;
  assign GEN_411 = 7'h9 == T_7300 ? T_7138_9 : GEN_410;
  assign GEN_412 = 7'ha == T_7300 ? T_7138_10 : GEN_411;
  assign GEN_413 = 7'hb == T_7300 ? T_7138_11 : GEN_412;
  assign GEN_414 = 7'hc == T_7300 ? T_7138_12 : GEN_413;
  assign GEN_415 = 7'hd == T_7300 ? T_7138_13 : GEN_414;
  assign GEN_416 = 7'he == T_7300 ? T_7138_14 : GEN_415;
  assign GEN_417 = 7'hf == T_7300 ? T_7138_15 : GEN_416;
  assign GEN_418 = 7'h10 == T_7300 ? T_7138_16 : GEN_417;
  assign GEN_419 = 7'h11 == T_7300 ? T_7138_17 : GEN_418;
  assign GEN_420 = 7'h12 == T_7300 ? T_7138_18 : GEN_419;
  assign GEN_421 = 7'h13 == T_7300 ? T_7138_19 : GEN_420;
  assign GEN_422 = 7'h14 == T_7300 ? T_7138_20 : GEN_421;
  assign GEN_423 = 7'h15 == T_7300 ? T_7138_21 : GEN_422;
  assign GEN_424 = 7'h16 == T_7300 ? T_7138_22 : GEN_423;
  assign GEN_425 = 7'h17 == T_7300 ? T_7138_23 : GEN_424;
  assign GEN_426 = 7'h18 == T_7300 ? T_7138_24 : GEN_425;
  assign GEN_427 = 7'h19 == T_7300 ? T_7138_25 : GEN_426;
  assign GEN_428 = 7'h1a == T_7300 ? T_7138_26 : GEN_427;
  assign GEN_429 = 7'h1b == T_7300 ? T_7138_27 : GEN_428;
  assign GEN_430 = 7'h1c == T_7300 ? T_7138_28 : GEN_429;
  assign GEN_431 = 7'h1d == T_7300 ? T_7138_29 : GEN_430;
  assign GEN_432 = 7'h1e == T_7300 ? T_7138_30 : GEN_431;
  assign GEN_433 = 7'h1f == T_7300 ? T_7138_31 : GEN_432;
  assign GEN_434 = 7'h20 == T_7300 ? T_7138_32 : GEN_433;
  assign GEN_435 = 7'h21 == T_7300 ? T_7138_33 : GEN_434;
  assign GEN_436 = 7'h22 == T_7300 ? T_7138_34 : GEN_435;
  assign GEN_437 = 7'h23 == T_7300 ? T_7138_35 : GEN_436;
  assign GEN_438 = 7'h24 == T_7300 ? T_7138_36 : GEN_437;
  assign GEN_439 = 7'h25 == T_7300 ? T_7138_37 : GEN_438;
  assign GEN_440 = 7'h26 == T_7300 ? T_7138_38 : GEN_439;
  assign GEN_441 = 7'h27 == T_7300 ? T_7138_39 : GEN_440;
  assign GEN_442 = 7'h28 == T_7300 ? T_7138_40 : GEN_441;
  assign GEN_443 = 7'h29 == T_7300 ? T_7138_41 : GEN_442;
  assign GEN_444 = 7'h2a == T_7300 ? T_7138_42 : GEN_443;
  assign GEN_445 = 7'h2b == T_7300 ? T_7138_43 : GEN_444;
  assign GEN_446 = 7'h2c == T_7300 ? T_7138_44 : GEN_445;
  assign GEN_447 = 7'h2d == T_7300 ? T_7138_45 : GEN_446;
  assign GEN_448 = 7'h2e == T_7300 ? T_7138_46 : GEN_447;
  assign GEN_449 = 7'h2f == T_7300 ? T_7138_47 : GEN_448;
  assign GEN_450 = 7'h30 == T_7300 ? T_7138_48 : GEN_449;
  assign GEN_451 = 7'h31 == T_7300 ? T_7138_49 : GEN_450;
  assign GEN_452 = 7'h32 == T_7300 ? T_7138_50 : GEN_451;
  assign GEN_453 = 7'h33 == T_7300 ? T_7138_51 : GEN_452;
  assign GEN_454 = 7'h34 == T_7300 ? T_7138_52 : GEN_453;
  assign GEN_455 = 7'h35 == T_7300 ? T_7138_53 : GEN_454;
  assign GEN_456 = 7'h36 == T_7300 ? T_7138_54 : GEN_455;
  assign GEN_457 = 7'h37 == T_7300 ? T_7138_55 : GEN_456;
  assign GEN_458 = 7'h38 == T_7300 ? T_7138_56 : GEN_457;
  assign GEN_459 = 7'h39 == T_7300 ? T_7138_57 : GEN_458;
  assign GEN_460 = 7'h3a == T_7300 ? T_7138_58 : GEN_459;
  assign GEN_461 = 7'h3b == T_7300 ? T_7138_59 : GEN_460;
  assign GEN_462 = 7'h3c == T_7300 ? T_7138_60 : GEN_461;
  assign GEN_463 = 7'h3d == T_7300 ? T_7138_61 : GEN_462;
  assign GEN_464 = 7'h3e == T_7300 ? T_7138_62 : GEN_463;
  assign GEN_465 = 7'h3f == T_7300 ? T_7138_63 : GEN_464;
  assign GEN_466 = 7'h40 == T_7300 ? T_7138_64 : GEN_465;
  assign GEN_467 = 7'h41 == T_7300 ? T_7138_65 : GEN_466;
  assign GEN_468 = 7'h42 == T_7300 ? T_7138_66 : GEN_467;
  assign GEN_469 = 7'h43 == T_7300 ? T_7138_67 : GEN_468;
  assign GEN_470 = 7'h44 == T_7300 ? T_7138_68 : GEN_469;
  assign GEN_471 = 7'h45 == T_7300 ? T_7138_69 : GEN_470;
  assign GEN_472 = 7'h46 == T_7300 ? T_7138_70 : GEN_471;
  assign GEN_473 = 7'h47 == T_7300 ? T_7138_71 : GEN_472;
  assign GEN_474 = 7'h48 == T_7300 ? T_7138_72 : GEN_473;
  assign GEN_475 = 7'h49 == T_7300 ? T_7138_73 : GEN_474;
  assign GEN_476 = 7'h4a == T_7300 ? T_7138_74 : GEN_475;
  assign GEN_477 = 7'h4b == T_7300 ? T_7138_75 : GEN_476;
  assign GEN_478 = 7'h4c == T_7300 ? T_7138_76 : GEN_477;
  assign GEN_479 = 7'h4d == T_7300 ? T_7138_77 : GEN_478;
  assign GEN_480 = 7'h4e == T_7300 ? T_7138_78 : GEN_479;
  assign GEN_481 = 7'h4f == T_7300 ? T_7138_79 : GEN_480;
  assign GEN_482 = 7'h50 == T_7300 ? T_7138_80 : GEN_481;
  assign GEN_483 = 7'h51 == T_7300 ? T_7138_81 : GEN_482;
  assign GEN_484 = 7'h52 == T_7300 ? T_7138_82 : GEN_483;
  assign GEN_485 = 7'h53 == T_7300 ? T_7138_83 : GEN_484;
  assign GEN_486 = 7'h54 == T_7300 ? T_7138_84 : GEN_485;
  assign GEN_487 = 7'h55 == T_7300 ? T_7138_85 : GEN_486;
  assign GEN_488 = 7'h56 == T_7300 ? T_7138_86 : GEN_487;
  assign GEN_489 = 7'h57 == T_7300 ? T_7138_87 : GEN_488;
  assign GEN_490 = 7'h58 == T_7300 ? T_7138_88 : GEN_489;
  assign GEN_491 = 7'h59 == T_7300 ? T_7138_89 : GEN_490;
  assign GEN_492 = 7'h5a == T_7300 ? T_7138_90 : GEN_491;
  assign GEN_493 = 7'h5b == T_7300 ? T_7138_91 : GEN_492;
  assign GEN_494 = 7'h5c == T_7300 ? T_7138_92 : GEN_493;
  assign GEN_495 = 7'h5d == T_7300 ? T_7138_93 : GEN_494;
  assign GEN_496 = 7'h5e == T_7300 ? T_7138_94 : GEN_495;
  assign GEN_497 = 7'h5f == T_7300 ? T_7138_95 : GEN_496;
  assign GEN_498 = 7'h60 == T_7300 ? T_7138_96 : GEN_497;
  assign GEN_499 = 7'h61 == T_7300 ? T_7138_97 : GEN_498;
  assign GEN_500 = 7'h62 == T_7300 ? T_7138_98 : GEN_499;
  assign GEN_501 = 7'h63 == T_7300 ? T_7138_99 : GEN_500;
  assign GEN_502 = 7'h64 == T_7300 ? T_7138_100 : GEN_501;
  assign GEN_503 = 7'h65 == T_7300 ? T_7138_101 : GEN_502;
  assign GEN_504 = 7'h66 == T_7300 ? T_7138_102 : GEN_503;
  assign GEN_505 = 7'h67 == T_7300 ? T_7138_103 : GEN_504;
  assign GEN_506 = 7'h68 == T_7300 ? T_7138_104 : GEN_505;
  assign GEN_507 = 7'h69 == T_7300 ? T_7138_105 : GEN_506;
  assign GEN_508 = 7'h6a == T_7300 ? T_7138_106 : GEN_507;
  assign GEN_509 = 7'h6b == T_7300 ? T_7138_107 : GEN_508;
  assign GEN_510 = 7'h6c == T_7300 ? T_7138_108 : GEN_509;
  assign GEN_511 = 7'h6d == T_7300 ? T_7138_109 : GEN_510;
  assign GEN_512 = 7'h6e == T_7300 ? T_7138_110 : GEN_511;
  assign GEN_513 = 7'h6f == T_7300 ? T_7138_111 : GEN_512;
  assign GEN_514 = 7'h70 == T_7300 ? T_7138_112 : GEN_513;
  assign GEN_515 = 7'h71 == T_7300 ? T_7138_113 : GEN_514;
  assign GEN_516 = 7'h72 == T_7300 ? T_7138_114 : GEN_515;
  assign GEN_517 = 7'h73 == T_7300 ? T_7138_115 : GEN_516;
  assign GEN_518 = 7'h74 == T_7300 ? T_7138_116 : GEN_517;
  assign GEN_519 = 7'h75 == T_7300 ? T_7138_117 : GEN_518;
  assign GEN_520 = 7'h76 == T_7300 ? T_7138_118 : GEN_519;
  assign GEN_521 = 7'h77 == T_7300 ? T_7138_119 : GEN_520;
  assign GEN_522 = 7'h78 == T_7300 ? T_7138_120 : GEN_521;
  assign GEN_523 = 7'h79 == T_7300 ? T_7138_121 : GEN_522;
  assign GEN_524 = 7'h7a == T_7300 ? T_7138_122 : GEN_523;
  assign GEN_525 = 7'h7b == T_7300 ? T_7138_123 : GEN_524;
  assign GEN_526 = 7'h7c == T_7300 ? T_7138_124 : GEN_525;
  assign GEN_527 = 7'h7d == T_7300 ? T_7138_125 : GEN_526;
  assign GEN_528 = 7'h7e == T_7300 ? T_7138_126 : GEN_527;
  assign GEN_529 = 7'h7f == T_7300 ? T_7138_127 : GEN_528;
  assign T_7306 = Queue_1_io_deq_bits_read ? GEN_2 : GEN_3;
  assign T_7307 = T_1028_ready & T_7303;
  assign T_7308 = T_953_valid & T_7303;
  assign T_7309 = T_992_ready & T_7306;
  assign T_7310 = Queue_1_io_deq_valid & T_7306;
  assign T_7312 = 128'h1 << T_7284;
  assign T_7313 = {1'h1,T_1322};
  assign T_7314 = {T_1583,T_1466};
  assign T_7315 = {T_7314,T_7313};
  assign T_7316 = {1'h1,T_1718};
  assign T_7317 = {T_1556,T_1394};
  assign T_7318 = {T_7317,T_7316};
  assign T_7319 = {T_7318,T_7315};
  assign T_7320 = {1'h1,T_1673};
  assign T_7322 = {2'h3,T_7320};
  assign T_7326 = {4'hf,T_7322};
  assign T_7327 = {T_7326,T_7319};
  assign T_7328 = {1'h1,T_1628};
  assign T_7329 = {T_1709,T_1610};
  assign T_7330 = {T_7329,T_7328};
  assign T_7331 = {1'h1,T_1358};
  assign T_7332 = {T_1664,T_1511};
  assign T_7333 = {T_7332,T_7331};
  assign T_7334 = {T_7333,T_7330};
  assign T_7335 = {1'h1,T_1340};
  assign T_7337 = {2'h3,T_7335};
  assign T_7341 = {4'hf,T_7337};
  assign T_7342 = {T_7341,T_7334};
  assign T_7343 = {T_7342,T_7327};
  assign T_7344 = {T_1421,T_1475};
  assign T_7345 = {T_1601,T_1484};
  assign T_7346 = {T_7345,T_7344};
  assign T_7347 = {T_1349,T_1700};
  assign T_7348 = {T_1565,T_1403};
  assign T_7349 = {T_7348,T_7347};
  assign T_7350 = {T_7349,T_7346};
  assign T_7351 = {T_1448,T_1655};
  assign T_7352 = {T_1646,T_1331};
  assign T_7353 = {T_7352,T_7351};
  assign T_7354 = {T_1493,T_1520};
  assign T_7355 = {T_1736,T_1367};
  assign T_7356 = {T_7355,T_7354};
  assign T_7357 = {T_7356,T_7353};
  assign T_7358 = {T_7357,T_7350};
  assign T_7374 = {16'hffff,T_7358};
  assign T_7375 = {T_7374,T_7343};
  assign T_7376 = {T_1430,T_1502};
  assign T_7377 = {T_1619,T_1574};
  assign T_7378 = {T_7377,T_7376};
  assign T_7379 = {T_1313,T_1745};
  assign T_7380 = {T_1529,T_1412};
  assign T_7381 = {T_7380,T_7379};
  assign T_7382 = {T_7381,T_7378};
  assign T_7383 = {T_1457,T_1637};
  assign T_7384 = {T_1682,T_1385};
  assign T_7385 = {T_7384,T_7383};
  assign T_7386 = {T_1439,T_1547};
  assign T_7387 = {T_1727,T_1376};
  assign T_7388 = {T_7387,T_7386};
  assign T_7389 = {T_7388,T_7385};
  assign T_7390 = {T_7389,T_7382};
  assign T_7391 = {T_1538,T_1592};
  assign T_7392 = {T_1754,T_1691};
  assign T_7393 = {T_7392,T_7391};
  assign T_7397 = {4'hf,T_7393};
  assign T_7405 = {8'hff,T_7397};
  assign T_7406 = {T_7405,T_7390};
  assign T_7438 = {32'hffffffff,T_7406};
  assign T_7439 = {T_7438,T_7375};
  assign T_7440 = T_7312 & T_7439;
  assign T_7442 = 128'h1 << T_7300;
  assign T_7443 = {1'h1,T_1326};
  assign T_7444 = {T_1587,T_1470};
  assign T_7445 = {T_7444,T_7443};
  assign T_7446 = {1'h1,T_1722};
  assign T_7447 = {T_1560,T_1398};
  assign T_7448 = {T_7447,T_7446};
  assign T_7449 = {T_7448,T_7445};
  assign T_7450 = {1'h1,T_1677};
  assign T_7452 = {2'h3,T_7450};
  assign T_7456 = {4'hf,T_7452};
  assign T_7457 = {T_7456,T_7449};
  assign T_7458 = {1'h1,T_1632};
  assign T_7459 = {T_1713,T_1614};
  assign T_7460 = {T_7459,T_7458};
  assign T_7461 = {1'h1,T_1362};
  assign T_7462 = {T_1668,T_1515};
  assign T_7463 = {T_7462,T_7461};
  assign T_7464 = {T_7463,T_7460};
  assign T_7465 = {1'h1,T_1344};
  assign T_7467 = {2'h3,T_7465};
  assign T_7471 = {4'hf,T_7467};
  assign T_7472 = {T_7471,T_7464};
  assign T_7473 = {T_7472,T_7457};
  assign T_7474 = {T_1425,T_1479};
  assign T_7475 = {T_1605,T_1488};
  assign T_7476 = {T_7475,T_7474};
  assign T_7477 = {T_1353,T_1704};
  assign T_7478 = {T_1569,T_1407};
  assign T_7479 = {T_7478,T_7477};
  assign T_7480 = {T_7479,T_7476};
  assign T_7481 = {T_1452,T_1659};
  assign T_7482 = {T_1650,T_1335};
  assign T_7483 = {T_7482,T_7481};
  assign T_7484 = {T_1497,T_1524};
  assign T_7485 = {T_1740,T_1371};
  assign T_7486 = {T_7485,T_7484};
  assign T_7487 = {T_7486,T_7483};
  assign T_7488 = {T_7487,T_7480};
  assign T_7504 = {16'hffff,T_7488};
  assign T_7505 = {T_7504,T_7473};
  assign T_7506 = {T_1434,T_1506};
  assign T_7507 = {T_1623,T_1578};
  assign T_7508 = {T_7507,T_7506};
  assign T_7509 = {T_1317,T_1749};
  assign T_7510 = {T_1533,T_1416};
  assign T_7511 = {T_7510,T_7509};
  assign T_7512 = {T_7511,T_7508};
  assign T_7513 = {T_1461,T_1641};
  assign T_7514 = {T_1686,T_1389};
  assign T_7515 = {T_7514,T_7513};
  assign T_7516 = {T_1443,T_1551};
  assign T_7517 = {T_1731,T_1380};
  assign T_7518 = {T_7517,T_7516};
  assign T_7519 = {T_7518,T_7515};
  assign T_7520 = {T_7519,T_7512};
  assign T_7521 = {T_1542,T_1596};
  assign T_7522 = {T_1758,T_1695};
  assign T_7523 = {T_7522,T_7521};
  assign T_7527 = {4'hf,T_7523};
  assign T_7535 = {8'hff,T_7527};
  assign T_7536 = {T_7535,T_7520};
  assign T_7568 = {32'hffffffff,T_7536};
  assign T_7569 = {T_7568,T_7505};
  assign T_7570 = T_7442 & T_7569;
  assign T_7571 = T_953_valid & T_1028_ready;
  assign T_7572 = T_7571 & T_1028_bits_read;
  assign T_7573 = T_7440[0];
  assign T_7574 = T_7572 & T_7573;
  assign T_7577 = T_1028_bits_read == 1'h0;
  assign T_7578 = T_7571 & T_7577;
  assign T_7580 = T_7578 & T_7573;
  assign T_7581 = Queue_1_io_deq_valid & T_992_ready;
  assign T_7582 = T_7581 & Queue_1_io_deq_bits_read;
  assign T_7583 = T_7570[0];
  assign T_7584 = T_7582 & T_7583;
  assign T_7587 = Queue_1_io_deq_bits_read == 1'h0;
  assign T_7588 = T_7581 & T_7587;
  assign T_7590 = T_7588 & T_7583;
  assign T_7613 = T_7440[2];
  assign T_7614 = T_7572 & T_7613;
  assign T_7620 = T_7578 & T_7613;
  assign T_7623 = T_7570[2];
  assign T_7624 = T_7582 & T_7623;
  assign T_7630 = T_7588 & T_7623;
  assign T_7633 = T_7440[3];
  assign T_7634 = T_7572 & T_7633;
  assign T_7640 = T_7578 & T_7633;
  assign T_7643 = T_7570[3];
  assign T_7644 = T_7582 & T_7643;
  assign T_7650 = T_7588 & T_7643;
  assign T_7653 = T_7440[4];
  assign T_7654 = T_7572 & T_7653;
  assign T_7660 = T_7578 & T_7653;
  assign T_7663 = T_7570[4];
  assign T_7664 = T_7582 & T_7663;
  assign T_7670 = T_7588 & T_7663;
  assign T_7693 = T_7440[6];
  assign T_7694 = T_7572 & T_7693;
  assign T_7700 = T_7578 & T_7693;
  assign T_7703 = T_7570[6];
  assign T_7704 = T_7582 & T_7703;
  assign T_7710 = T_7588 & T_7703;
  assign T_7713 = T_7440[7];
  assign T_7714 = T_7572 & T_7713;
  assign T_7720 = T_7578 & T_7713;
  assign T_7723 = T_7570[7];
  assign T_7724 = T_7582 & T_7723;
  assign T_7730 = T_7588 & T_7723;
  assign T_7733 = T_7440[8];
  assign T_7734 = T_7572 & T_7733;
  assign T_7740 = T_7578 & T_7733;
  assign T_7743 = T_7570[8];
  assign T_7744 = T_7582 & T_7743;
  assign T_7750 = T_7588 & T_7743;
  assign T_7893 = T_7440[16];
  assign T_7894 = T_7572 & T_7893;
  assign T_7900 = T_7578 & T_7893;
  assign T_7903 = T_7570[16];
  assign T_7904 = T_7582 & T_7903;
  assign T_7910 = T_7588 & T_7903;
  assign T_7933 = T_7440[18];
  assign T_7934 = T_7572 & T_7933;
  assign T_7940 = T_7578 & T_7933;
  assign T_7943 = T_7570[18];
  assign T_7944 = T_7582 & T_7943;
  assign T_7950 = T_7588 & T_7943;
  assign T_7953 = T_7440[19];
  assign T_7954 = T_7572 & T_7953;
  assign T_7960 = T_7578 & T_7953;
  assign T_7963 = T_7570[19];
  assign T_7964 = T_7582 & T_7963;
  assign T_7970 = T_7588 & T_7963;
  assign T_7973 = T_7440[20];
  assign T_7974 = T_7572 & T_7973;
  assign T_7980 = T_7578 & T_7973;
  assign T_7983 = T_7570[20];
  assign T_7984 = T_7582 & T_7983;
  assign T_7990 = T_7588 & T_7983;
  assign T_8013 = T_7440[22];
  assign T_8014 = T_7572 & T_8013;
  assign T_8020 = T_7578 & T_8013;
  assign T_8023 = T_7570[22];
  assign T_8024 = T_7582 & T_8023;
  assign T_8030 = T_7588 & T_8023;
  assign T_8033 = T_7440[23];
  assign T_8034 = T_7572 & T_8033;
  assign T_8040 = T_7578 & T_8033;
  assign T_8043 = T_7570[23];
  assign T_8044 = T_7582 & T_8043;
  assign T_8050 = T_7588 & T_8043;
  assign T_8053 = T_7440[24];
  assign T_8054 = T_7572 & T_8053;
  assign T_8060 = T_7578 & T_8053;
  assign T_8063 = T_7570[24];
  assign T_8064 = T_7582 & T_8063;
  assign T_8070 = T_7588 & T_8063;
  assign T_8213 = T_7440[32];
  assign T_8214 = T_7572 & T_8213;
  assign T_8220 = T_7578 & T_8213;
  assign T_8223 = T_7570[32];
  assign T_8224 = T_7582 & T_8223;
  assign T_8230 = T_7588 & T_8223;
  assign T_8233 = T_7440[33];
  assign T_8234 = T_7572 & T_8233;
  assign T_8240 = T_7578 & T_8233;
  assign T_8243 = T_7570[33];
  assign T_8244 = T_7582 & T_8243;
  assign T_8250 = T_7588 & T_8243;
  assign T_8253 = T_7440[34];
  assign T_8254 = T_7572 & T_8253;
  assign T_8260 = T_7578 & T_8253;
  assign T_8263 = T_7570[34];
  assign T_8264 = T_7582 & T_8263;
  assign T_8270 = T_7588 & T_8263;
  assign T_8273 = T_7440[35];
  assign T_8274 = T_7572 & T_8273;
  assign T_8280 = T_7578 & T_8273;
  assign T_8283 = T_7570[35];
  assign T_8284 = T_7582 & T_8283;
  assign T_8290 = T_7588 & T_8283;
  assign T_8293 = T_7440[36];
  assign T_8294 = T_7572 & T_8293;
  assign T_8300 = T_7578 & T_8293;
  assign T_8303 = T_7570[36];
  assign T_8304 = T_7582 & T_8303;
  assign T_8310 = T_7588 & T_8303;
  assign T_8313 = T_7440[37];
  assign T_8314 = T_7572 & T_8313;
  assign T_8320 = T_7578 & T_8313;
  assign T_8323 = T_7570[37];
  assign T_8324 = T_7582 & T_8323;
  assign T_8330 = T_7588 & T_8323;
  assign T_8333 = T_7440[38];
  assign T_8334 = T_7572 & T_8333;
  assign T_8340 = T_7578 & T_8333;
  assign T_8343 = T_7570[38];
  assign T_8344 = T_7582 & T_8343;
  assign T_8350 = T_7588 & T_8343;
  assign T_8353 = T_7440[39];
  assign T_8354 = T_7572 & T_8353;
  assign T_8360 = T_7578 & T_8353;
  assign T_8363 = T_7570[39];
  assign T_8364 = T_7582 & T_8363;
  assign T_8370 = T_7588 & T_8363;
  assign T_8373 = T_7440[40];
  assign T_8374 = T_7572 & T_8373;
  assign T_8380 = T_7578 & T_8373;
  assign T_8383 = T_7570[40];
  assign T_8384 = T_7582 & T_8383;
  assign T_8390 = T_7588 & T_8383;
  assign T_8393 = T_7440[41];
  assign T_8394 = T_7572 & T_8393;
  assign T_8400 = T_7578 & T_8393;
  assign T_8403 = T_7570[41];
  assign T_8404 = T_7582 & T_8403;
  assign T_8410 = T_7588 & T_8403;
  assign T_8413 = T_7440[42];
  assign T_8414 = T_7572 & T_8413;
  assign T_8420 = T_7578 & T_8413;
  assign T_8423 = T_7570[42];
  assign T_8424 = T_7582 & T_8423;
  assign T_8430 = T_7588 & T_8423;
  assign T_8433 = T_7440[43];
  assign T_8434 = T_7572 & T_8433;
  assign T_8440 = T_7578 & T_8433;
  assign T_8443 = T_7570[43];
  assign T_8444 = T_7582 & T_8443;
  assign T_8450 = T_7588 & T_8443;
  assign T_8453 = T_7440[44];
  assign T_8454 = T_7572 & T_8453;
  assign T_8460 = T_7578 & T_8453;
  assign T_8463 = T_7570[44];
  assign T_8464 = T_7582 & T_8463;
  assign T_8470 = T_7588 & T_8463;
  assign T_8473 = T_7440[45];
  assign T_8474 = T_7572 & T_8473;
  assign T_8480 = T_7578 & T_8473;
  assign T_8483 = T_7570[45];
  assign T_8484 = T_7582 & T_8483;
  assign T_8490 = T_7588 & T_8483;
  assign T_8493 = T_7440[46];
  assign T_8494 = T_7572 & T_8493;
  assign T_8500 = T_7578 & T_8493;
  assign T_8503 = T_7570[46];
  assign T_8504 = T_7582 & T_8503;
  assign T_8510 = T_7588 & T_8503;
  assign T_8513 = T_7440[47];
  assign T_8514 = T_7572 & T_8513;
  assign T_8520 = T_7578 & T_8513;
  assign T_8523 = T_7570[47];
  assign T_8524 = T_7582 & T_8523;
  assign T_8530 = T_7588 & T_8523;
  assign T_8853 = T_7440[64];
  assign T_8854 = T_7572 & T_8853;
  assign T_8860 = T_7578 & T_8853;
  assign T_8863 = T_7570[64];
  assign T_8864 = T_7582 & T_8863;
  assign T_8870 = T_7588 & T_8863;
  assign T_8873 = T_7440[65];
  assign T_8874 = T_7572 & T_8873;
  assign T_8880 = T_7578 & T_8873;
  assign T_8883 = T_7570[65];
  assign T_8884 = T_7582 & T_8883;
  assign T_8890 = T_7588 & T_8883;
  assign T_8893 = T_7440[66];
  assign T_8894 = T_7572 & T_8893;
  assign T_8900 = T_7578 & T_8893;
  assign T_8903 = T_7570[66];
  assign T_8904 = T_7582 & T_8903;
  assign T_8910 = T_7588 & T_8903;
  assign T_8913 = T_7440[67];
  assign T_8914 = T_7572 & T_8913;
  assign T_8920 = T_7578 & T_8913;
  assign T_8923 = T_7570[67];
  assign T_8924 = T_7582 & T_8923;
  assign T_8930 = T_7588 & T_8923;
  assign T_8933 = T_7440[68];
  assign T_8934 = T_7572 & T_8933;
  assign T_8940 = T_7578 & T_8933;
  assign T_8943 = T_7570[68];
  assign T_8944 = T_7582 & T_8943;
  assign T_8950 = T_7588 & T_8943;
  assign T_8953 = T_7440[69];
  assign T_8954 = T_7572 & T_8953;
  assign T_8960 = T_7578 & T_8953;
  assign T_8963 = T_7570[69];
  assign T_8964 = T_7582 & T_8963;
  assign T_8970 = T_7588 & T_8963;
  assign T_8973 = T_7440[70];
  assign T_8974 = T_7572 & T_8973;
  assign T_8980 = T_7578 & T_8973;
  assign T_8983 = T_7570[70];
  assign T_8984 = T_7582 & T_8983;
  assign T_8990 = T_7588 & T_8983;
  assign T_8993 = T_7440[71];
  assign T_8994 = T_7572 & T_8993;
  assign T_9000 = T_7578 & T_8993;
  assign T_9003 = T_7570[71];
  assign T_9004 = T_7582 & T_9003;
  assign T_9010 = T_7588 & T_9003;
  assign T_9013 = T_7440[72];
  assign T_9014 = T_7572 & T_9013;
  assign T_9020 = T_7578 & T_9013;
  assign T_9023 = T_7570[72];
  assign T_9024 = T_7582 & T_9023;
  assign T_9030 = T_7588 & T_9023;
  assign T_9033 = T_7440[73];
  assign T_9034 = T_7572 & T_9033;
  assign T_9040 = T_7578 & T_9033;
  assign T_9043 = T_7570[73];
  assign T_9044 = T_7582 & T_9043;
  assign T_9050 = T_7588 & T_9043;
  assign T_9053 = T_7440[74];
  assign T_9054 = T_7572 & T_9053;
  assign T_9060 = T_7578 & T_9053;
  assign T_9063 = T_7570[74];
  assign T_9064 = T_7582 & T_9063;
  assign T_9070 = T_7588 & T_9063;
  assign T_9073 = T_7440[75];
  assign T_9074 = T_7572 & T_9073;
  assign T_9080 = T_7578 & T_9073;
  assign T_9083 = T_7570[75];
  assign T_9084 = T_7582 & T_9083;
  assign T_9090 = T_7588 & T_9083;
  assign T_9093 = T_7440[76];
  assign T_9094 = T_7572 & T_9093;
  assign T_9100 = T_7578 & T_9093;
  assign T_9103 = T_7570[76];
  assign T_9104 = T_7582 & T_9103;
  assign T_9110 = T_7588 & T_9103;
  assign T_9113 = T_7440[77];
  assign T_9114 = T_7572 & T_9113;
  assign T_9120 = T_7578 & T_9113;
  assign T_9123 = T_7570[77];
  assign T_9124 = T_7582 & T_9123;
  assign T_9130 = T_7588 & T_9123;
  assign T_9133 = T_7440[78];
  assign T_9134 = T_7572 & T_9133;
  assign T_9140 = T_7578 & T_9133;
  assign T_9143 = T_7570[78];
  assign T_9144 = T_7582 & T_9143;
  assign T_9150 = T_7588 & T_9143;
  assign T_9153 = T_7440[79];
  assign T_9154 = T_7572 & T_9153;
  assign T_9160 = T_7578 & T_9153;
  assign T_9163 = T_7570[79];
  assign T_9164 = T_7582 & T_9163;
  assign T_9170 = T_7588 & T_9163;
  assign T_9173 = T_7440[80];
  assign T_9174 = T_7572 & T_9173;
  assign T_9180 = T_7578 & T_9173;
  assign T_9183 = T_7570[80];
  assign T_9184 = T_7582 & T_9183;
  assign T_9190 = T_7588 & T_9183;
  assign T_9193 = T_7440[81];
  assign T_9194 = T_7572 & T_9193;
  assign T_9200 = T_7578 & T_9193;
  assign T_9203 = T_7570[81];
  assign T_9204 = T_7582 & T_9203;
  assign T_9210 = T_7588 & T_9203;
  assign T_9213 = T_7440[82];
  assign T_9214 = T_7572 & T_9213;
  assign T_9220 = T_7578 & T_9213;
  assign T_9223 = T_7570[82];
  assign T_9224 = T_7582 & T_9223;
  assign T_9230 = T_7588 & T_9223;
  assign T_9233 = T_7440[83];
  assign T_9234 = T_7572 & T_9233;
  assign T_9240 = T_7578 & T_9233;
  assign T_9243 = T_7570[83];
  assign T_9244 = T_7582 & T_9243;
  assign T_9250 = T_7588 & T_9243;
  assign T_10462_0 = T_1326;
  assign T_10462_1 = 1'h1;
  assign T_10462_2 = T_1470;
  assign T_10462_3 = T_1587;
  assign T_10462_4 = T_1722;
  assign T_10462_5 = 1'h1;
  assign T_10462_6 = T_1398;
  assign T_10462_7 = T_1560;
  assign T_10462_8 = T_1677;
  assign T_10462_9 = 1'h1;
  assign T_10462_10 = 1'h1;
  assign T_10462_11 = 1'h1;
  assign T_10462_12 = 1'h1;
  assign T_10462_13 = 1'h1;
  assign T_10462_14 = 1'h1;
  assign T_10462_15 = 1'h1;
  assign T_10462_16 = T_1632;
  assign T_10462_17 = 1'h1;
  assign T_10462_18 = T_1614;
  assign T_10462_19 = T_1713;
  assign T_10462_20 = T_1362;
  assign T_10462_21 = 1'h1;
  assign T_10462_22 = T_1515;
  assign T_10462_23 = T_1668;
  assign T_10462_24 = T_1344;
  assign T_10462_25 = 1'h1;
  assign T_10462_26 = 1'h1;
  assign T_10462_27 = 1'h1;
  assign T_10462_28 = 1'h1;
  assign T_10462_29 = 1'h1;
  assign T_10462_30 = 1'h1;
  assign T_10462_31 = 1'h1;
  assign T_10462_32 = T_1479;
  assign T_10462_33 = T_1425;
  assign T_10462_34 = T_1488;
  assign T_10462_35 = T_1605;
  assign T_10462_36 = T_1704;
  assign T_10462_37 = T_1353;
  assign T_10462_38 = T_1407;
  assign T_10462_39 = T_1569;
  assign T_10462_40 = T_1659;
  assign T_10462_41 = T_1452;
  assign T_10462_42 = T_1335;
  assign T_10462_43 = T_1650;
  assign T_10462_44 = T_1524;
  assign T_10462_45 = T_1497;
  assign T_10462_46 = T_1371;
  assign T_10462_47 = T_1740;
  assign T_10462_48 = 1'h1;
  assign T_10462_49 = 1'h1;
  assign T_10462_50 = 1'h1;
  assign T_10462_51 = 1'h1;
  assign T_10462_52 = 1'h1;
  assign T_10462_53 = 1'h1;
  assign T_10462_54 = 1'h1;
  assign T_10462_55 = 1'h1;
  assign T_10462_56 = 1'h1;
  assign T_10462_57 = 1'h1;
  assign T_10462_58 = 1'h1;
  assign T_10462_59 = 1'h1;
  assign T_10462_60 = 1'h1;
  assign T_10462_61 = 1'h1;
  assign T_10462_62 = 1'h1;
  assign T_10462_63 = 1'h1;
  assign T_10462_64 = T_1506;
  assign T_10462_65 = T_1434;
  assign T_10462_66 = T_1578;
  assign T_10462_67 = T_1623;
  assign T_10462_68 = T_1749;
  assign T_10462_69 = T_1317;
  assign T_10462_70 = T_1416;
  assign T_10462_71 = T_1533;
  assign T_10462_72 = T_1641;
  assign T_10462_73 = T_1461;
  assign T_10462_74 = T_1389;
  assign T_10462_75 = T_1686;
  assign T_10462_76 = T_1551;
  assign T_10462_77 = T_1443;
  assign T_10462_78 = T_1380;
  assign T_10462_79 = T_1731;
  assign T_10462_80 = T_1596;
  assign T_10462_81 = T_1542;
  assign T_10462_82 = T_1695;
  assign T_10462_83 = T_1758;
  assign T_10462_84 = 1'h1;
  assign T_10462_85 = 1'h1;
  assign T_10462_86 = 1'h1;
  assign T_10462_87 = 1'h1;
  assign T_10462_88 = 1'h1;
  assign T_10462_89 = 1'h1;
  assign T_10462_90 = 1'h1;
  assign T_10462_91 = 1'h1;
  assign T_10462_92 = 1'h1;
  assign T_10462_93 = 1'h1;
  assign T_10462_94 = 1'h1;
  assign T_10462_95 = 1'h1;
  assign T_10462_96 = 1'h1;
  assign T_10462_97 = 1'h1;
  assign T_10462_98 = 1'h1;
  assign T_10462_99 = 1'h1;
  assign T_10462_100 = 1'h1;
  assign T_10462_101 = 1'h1;
  assign T_10462_102 = 1'h1;
  assign T_10462_103 = 1'h1;
  assign T_10462_104 = 1'h1;
  assign T_10462_105 = 1'h1;
  assign T_10462_106 = 1'h1;
  assign T_10462_107 = 1'h1;
  assign T_10462_108 = 1'h1;
  assign T_10462_109 = 1'h1;
  assign T_10462_110 = 1'h1;
  assign T_10462_111 = 1'h1;
  assign T_10462_112 = 1'h1;
  assign T_10462_113 = 1'h1;
  assign T_10462_114 = 1'h1;
  assign T_10462_115 = 1'h1;
  assign T_10462_116 = 1'h1;
  assign T_10462_117 = 1'h1;
  assign T_10462_118 = 1'h1;
  assign T_10462_119 = 1'h1;
  assign T_10462_120 = 1'h1;
  assign T_10462_121 = 1'h1;
  assign T_10462_122 = 1'h1;
  assign T_10462_123 = 1'h1;
  assign T_10462_124 = 1'h1;
  assign T_10462_125 = 1'h1;
  assign T_10462_126 = 1'h1;
  assign T_10462_127 = 1'h1;
  assign T_10725_0 = T_2560;
  assign T_10725_1 = 32'h0;
  assign T_10725_2 = T_3200;
  assign T_10725_3 = T_3720;
  assign T_10725_4 = {{16'd0}, T_4320};
  assign T_10725_5 = 32'h0;
  assign T_10725_6 = T_2880;
  assign T_10725_7 = T_3600;
  assign T_10725_8 = {{16'd0}, T_4120};
  assign T_10725_9 = 32'h0;
  assign T_10725_10 = 32'h0;
  assign T_10725_11 = 32'h0;
  assign T_10725_12 = 32'h0;
  assign T_10725_13 = 32'h0;
  assign T_10725_14 = 32'h0;
  assign T_10725_15 = 32'h0;
  assign T_10725_16 = T_3920;
  assign T_10725_17 = 32'h0;
  assign T_10725_18 = T_3840;
  assign T_10725_19 = T_4280;
  assign T_10725_20 = T_2720;
  assign T_10725_21 = 32'h0;
  assign T_10725_22 = T_3400;
  assign T_10725_23 = T_4080;
  assign T_10725_24 = T_2640;
  assign T_10725_25 = 32'h0;
  assign T_10725_26 = 32'h0;
  assign T_10725_27 = 32'h0;
  assign T_10725_28 = 32'h0;
  assign T_10725_29 = 32'h0;
  assign T_10725_30 = 32'h0;
  assign T_10725_31 = 32'h0;
  assign T_10725_32 = backupRegs_0;
  assign T_10725_33 = backupRegs_1;
  assign T_10725_34 = backupRegs_2;
  assign T_10725_35 = backupRegs_3;
  assign T_10725_36 = backupRegs_4;
  assign T_10725_37 = backupRegs_5;
  assign T_10725_38 = backupRegs_6;
  assign T_10725_39 = backupRegs_7;
  assign T_10725_40 = backupRegs_8;
  assign T_10725_41 = backupRegs_9;
  assign T_10725_42 = backupRegs_10;
  assign T_10725_43 = backupRegs_11;
  assign T_10725_44 = backupRegs_12;
  assign T_10725_45 = backupRegs_13;
  assign T_10725_46 = backupRegs_14;
  assign T_10725_47 = backupRegs_15;
  assign T_10725_48 = 32'h0;
  assign T_10725_49 = 32'h0;
  assign T_10725_50 = 32'h0;
  assign T_10725_51 = 32'h0;
  assign T_10725_52 = 32'h0;
  assign T_10725_53 = 32'h0;
  assign T_10725_54 = 32'h0;
  assign T_10725_55 = 32'h0;
  assign T_10725_56 = 32'h0;
  assign T_10725_57 = 32'h0;
  assign T_10725_58 = 32'h0;
  assign T_10725_59 = 32'h0;
  assign T_10725_60 = 32'h0;
  assign T_10725_61 = 32'h0;
  assign T_10725_62 = 32'h0;
  assign T_10725_63 = 32'h0;
  assign T_10725_64 = T_3360;
  assign T_10725_65 = T_3040;
  assign T_10725_66 = T_3680;
  assign T_10725_67 = T_3880;
  assign T_10725_68 = T_4440;
  assign T_10725_69 = T_2520;
  assign T_10725_70 = T_2960;
  assign T_10725_71 = T_3480;
  assign T_10725_72 = T_3960;
  assign T_10725_73 = T_3160;
  assign T_10725_74 = T_2840;
  assign T_10725_75 = T_4160;
  assign T_10725_76 = T_3560;
  assign T_10725_77 = T_3080;
  assign T_10725_78 = T_2800;
  assign T_10725_79 = T_4360;
  assign T_10725_80 = {{28'd0}, T_3760};
  assign T_10725_81 = T_3520;
  assign T_10725_82 = T_4200;
  assign T_10725_83 = T_4480;
  assign T_10725_84 = 32'h0;
  assign T_10725_85 = 32'h0;
  assign T_10725_86 = 32'h0;
  assign T_10725_87 = 32'h0;
  assign T_10725_88 = 32'h0;
  assign T_10725_89 = 32'h0;
  assign T_10725_90 = 32'h0;
  assign T_10725_91 = 32'h0;
  assign T_10725_92 = 32'h0;
  assign T_10725_93 = 32'h0;
  assign T_10725_94 = 32'h0;
  assign T_10725_95 = 32'h0;
  assign T_10725_96 = 32'h0;
  assign T_10725_97 = 32'h0;
  assign T_10725_98 = 32'h0;
  assign T_10725_99 = 32'h0;
  assign T_10725_100 = 32'h0;
  assign T_10725_101 = 32'h0;
  assign T_10725_102 = 32'h0;
  assign T_10725_103 = 32'h0;
  assign T_10725_104 = 32'h0;
  assign T_10725_105 = 32'h0;
  assign T_10725_106 = 32'h0;
  assign T_10725_107 = 32'h0;
  assign T_10725_108 = 32'h0;
  assign T_10725_109 = 32'h0;
  assign T_10725_110 = 32'h0;
  assign T_10725_111 = 32'h0;
  assign T_10725_112 = 32'h0;
  assign T_10725_113 = 32'h0;
  assign T_10725_114 = 32'h0;
  assign T_10725_115 = 32'h0;
  assign T_10725_116 = 32'h0;
  assign T_10725_117 = 32'h0;
  assign T_10725_118 = 32'h0;
  assign T_10725_119 = 32'h0;
  assign T_10725_120 = 32'h0;
  assign T_10725_121 = 32'h0;
  assign T_10725_122 = 32'h0;
  assign T_10725_123 = 32'h0;
  assign T_10725_124 = 32'h0;
  assign T_10725_125 = 32'h0;
  assign T_10725_126 = 32'h0;
  assign T_10725_127 = 32'h0;
  assign GEN_4 = GEN_656;
  assign GEN_530 = 7'h1 == T_7300 ? T_10462_1 : T_10462_0;
  assign GEN_531 = 7'h2 == T_7300 ? T_10462_2 : GEN_530;
  assign GEN_532 = 7'h3 == T_7300 ? T_10462_3 : GEN_531;
  assign GEN_533 = 7'h4 == T_7300 ? T_10462_4 : GEN_532;
  assign GEN_534 = 7'h5 == T_7300 ? T_10462_5 : GEN_533;
  assign GEN_535 = 7'h6 == T_7300 ? T_10462_6 : GEN_534;
  assign GEN_536 = 7'h7 == T_7300 ? T_10462_7 : GEN_535;
  assign GEN_537 = 7'h8 == T_7300 ? T_10462_8 : GEN_536;
  assign GEN_538 = 7'h9 == T_7300 ? T_10462_9 : GEN_537;
  assign GEN_539 = 7'ha == T_7300 ? T_10462_10 : GEN_538;
  assign GEN_540 = 7'hb == T_7300 ? T_10462_11 : GEN_539;
  assign GEN_541 = 7'hc == T_7300 ? T_10462_12 : GEN_540;
  assign GEN_542 = 7'hd == T_7300 ? T_10462_13 : GEN_541;
  assign GEN_543 = 7'he == T_7300 ? T_10462_14 : GEN_542;
  assign GEN_544 = 7'hf == T_7300 ? T_10462_15 : GEN_543;
  assign GEN_545 = 7'h10 == T_7300 ? T_10462_16 : GEN_544;
  assign GEN_546 = 7'h11 == T_7300 ? T_10462_17 : GEN_545;
  assign GEN_547 = 7'h12 == T_7300 ? T_10462_18 : GEN_546;
  assign GEN_548 = 7'h13 == T_7300 ? T_10462_19 : GEN_547;
  assign GEN_549 = 7'h14 == T_7300 ? T_10462_20 : GEN_548;
  assign GEN_550 = 7'h15 == T_7300 ? T_10462_21 : GEN_549;
  assign GEN_551 = 7'h16 == T_7300 ? T_10462_22 : GEN_550;
  assign GEN_552 = 7'h17 == T_7300 ? T_10462_23 : GEN_551;
  assign GEN_553 = 7'h18 == T_7300 ? T_10462_24 : GEN_552;
  assign GEN_554 = 7'h19 == T_7300 ? T_10462_25 : GEN_553;
  assign GEN_555 = 7'h1a == T_7300 ? T_10462_26 : GEN_554;
  assign GEN_556 = 7'h1b == T_7300 ? T_10462_27 : GEN_555;
  assign GEN_557 = 7'h1c == T_7300 ? T_10462_28 : GEN_556;
  assign GEN_558 = 7'h1d == T_7300 ? T_10462_29 : GEN_557;
  assign GEN_559 = 7'h1e == T_7300 ? T_10462_30 : GEN_558;
  assign GEN_560 = 7'h1f == T_7300 ? T_10462_31 : GEN_559;
  assign GEN_561 = 7'h20 == T_7300 ? T_10462_32 : GEN_560;
  assign GEN_562 = 7'h21 == T_7300 ? T_10462_33 : GEN_561;
  assign GEN_563 = 7'h22 == T_7300 ? T_10462_34 : GEN_562;
  assign GEN_564 = 7'h23 == T_7300 ? T_10462_35 : GEN_563;
  assign GEN_565 = 7'h24 == T_7300 ? T_10462_36 : GEN_564;
  assign GEN_566 = 7'h25 == T_7300 ? T_10462_37 : GEN_565;
  assign GEN_567 = 7'h26 == T_7300 ? T_10462_38 : GEN_566;
  assign GEN_568 = 7'h27 == T_7300 ? T_10462_39 : GEN_567;
  assign GEN_569 = 7'h28 == T_7300 ? T_10462_40 : GEN_568;
  assign GEN_570 = 7'h29 == T_7300 ? T_10462_41 : GEN_569;
  assign GEN_571 = 7'h2a == T_7300 ? T_10462_42 : GEN_570;
  assign GEN_572 = 7'h2b == T_7300 ? T_10462_43 : GEN_571;
  assign GEN_573 = 7'h2c == T_7300 ? T_10462_44 : GEN_572;
  assign GEN_574 = 7'h2d == T_7300 ? T_10462_45 : GEN_573;
  assign GEN_575 = 7'h2e == T_7300 ? T_10462_46 : GEN_574;
  assign GEN_576 = 7'h2f == T_7300 ? T_10462_47 : GEN_575;
  assign GEN_577 = 7'h30 == T_7300 ? T_10462_48 : GEN_576;
  assign GEN_578 = 7'h31 == T_7300 ? T_10462_49 : GEN_577;
  assign GEN_579 = 7'h32 == T_7300 ? T_10462_50 : GEN_578;
  assign GEN_580 = 7'h33 == T_7300 ? T_10462_51 : GEN_579;
  assign GEN_581 = 7'h34 == T_7300 ? T_10462_52 : GEN_580;
  assign GEN_582 = 7'h35 == T_7300 ? T_10462_53 : GEN_581;
  assign GEN_583 = 7'h36 == T_7300 ? T_10462_54 : GEN_582;
  assign GEN_584 = 7'h37 == T_7300 ? T_10462_55 : GEN_583;
  assign GEN_585 = 7'h38 == T_7300 ? T_10462_56 : GEN_584;
  assign GEN_586 = 7'h39 == T_7300 ? T_10462_57 : GEN_585;
  assign GEN_587 = 7'h3a == T_7300 ? T_10462_58 : GEN_586;
  assign GEN_588 = 7'h3b == T_7300 ? T_10462_59 : GEN_587;
  assign GEN_589 = 7'h3c == T_7300 ? T_10462_60 : GEN_588;
  assign GEN_590 = 7'h3d == T_7300 ? T_10462_61 : GEN_589;
  assign GEN_591 = 7'h3e == T_7300 ? T_10462_62 : GEN_590;
  assign GEN_592 = 7'h3f == T_7300 ? T_10462_63 : GEN_591;
  assign GEN_593 = 7'h40 == T_7300 ? T_10462_64 : GEN_592;
  assign GEN_594 = 7'h41 == T_7300 ? T_10462_65 : GEN_593;
  assign GEN_595 = 7'h42 == T_7300 ? T_10462_66 : GEN_594;
  assign GEN_596 = 7'h43 == T_7300 ? T_10462_67 : GEN_595;
  assign GEN_597 = 7'h44 == T_7300 ? T_10462_68 : GEN_596;
  assign GEN_598 = 7'h45 == T_7300 ? T_10462_69 : GEN_597;
  assign GEN_599 = 7'h46 == T_7300 ? T_10462_70 : GEN_598;
  assign GEN_600 = 7'h47 == T_7300 ? T_10462_71 : GEN_599;
  assign GEN_601 = 7'h48 == T_7300 ? T_10462_72 : GEN_600;
  assign GEN_602 = 7'h49 == T_7300 ? T_10462_73 : GEN_601;
  assign GEN_603 = 7'h4a == T_7300 ? T_10462_74 : GEN_602;
  assign GEN_604 = 7'h4b == T_7300 ? T_10462_75 : GEN_603;
  assign GEN_605 = 7'h4c == T_7300 ? T_10462_76 : GEN_604;
  assign GEN_606 = 7'h4d == T_7300 ? T_10462_77 : GEN_605;
  assign GEN_607 = 7'h4e == T_7300 ? T_10462_78 : GEN_606;
  assign GEN_608 = 7'h4f == T_7300 ? T_10462_79 : GEN_607;
  assign GEN_609 = 7'h50 == T_7300 ? T_10462_80 : GEN_608;
  assign GEN_610 = 7'h51 == T_7300 ? T_10462_81 : GEN_609;
  assign GEN_611 = 7'h52 == T_7300 ? T_10462_82 : GEN_610;
  assign GEN_612 = 7'h53 == T_7300 ? T_10462_83 : GEN_611;
  assign GEN_613 = 7'h54 == T_7300 ? T_10462_84 : GEN_612;
  assign GEN_614 = 7'h55 == T_7300 ? T_10462_85 : GEN_613;
  assign GEN_615 = 7'h56 == T_7300 ? T_10462_86 : GEN_614;
  assign GEN_616 = 7'h57 == T_7300 ? T_10462_87 : GEN_615;
  assign GEN_617 = 7'h58 == T_7300 ? T_10462_88 : GEN_616;
  assign GEN_618 = 7'h59 == T_7300 ? T_10462_89 : GEN_617;
  assign GEN_619 = 7'h5a == T_7300 ? T_10462_90 : GEN_618;
  assign GEN_620 = 7'h5b == T_7300 ? T_10462_91 : GEN_619;
  assign GEN_621 = 7'h5c == T_7300 ? T_10462_92 : GEN_620;
  assign GEN_622 = 7'h5d == T_7300 ? T_10462_93 : GEN_621;
  assign GEN_623 = 7'h5e == T_7300 ? T_10462_94 : GEN_622;
  assign GEN_624 = 7'h5f == T_7300 ? T_10462_95 : GEN_623;
  assign GEN_625 = 7'h60 == T_7300 ? T_10462_96 : GEN_624;
  assign GEN_626 = 7'h61 == T_7300 ? T_10462_97 : GEN_625;
  assign GEN_627 = 7'h62 == T_7300 ? T_10462_98 : GEN_626;
  assign GEN_628 = 7'h63 == T_7300 ? T_10462_99 : GEN_627;
  assign GEN_629 = 7'h64 == T_7300 ? T_10462_100 : GEN_628;
  assign GEN_630 = 7'h65 == T_7300 ? T_10462_101 : GEN_629;
  assign GEN_631 = 7'h66 == T_7300 ? T_10462_102 : GEN_630;
  assign GEN_632 = 7'h67 == T_7300 ? T_10462_103 : GEN_631;
  assign GEN_633 = 7'h68 == T_7300 ? T_10462_104 : GEN_632;
  assign GEN_634 = 7'h69 == T_7300 ? T_10462_105 : GEN_633;
  assign GEN_635 = 7'h6a == T_7300 ? T_10462_106 : GEN_634;
  assign GEN_636 = 7'h6b == T_7300 ? T_10462_107 : GEN_635;
  assign GEN_637 = 7'h6c == T_7300 ? T_10462_108 : GEN_636;
  assign GEN_638 = 7'h6d == T_7300 ? T_10462_109 : GEN_637;
  assign GEN_639 = 7'h6e == T_7300 ? T_10462_110 : GEN_638;
  assign GEN_640 = 7'h6f == T_7300 ? T_10462_111 : GEN_639;
  assign GEN_641 = 7'h70 == T_7300 ? T_10462_112 : GEN_640;
  assign GEN_642 = 7'h71 == T_7300 ? T_10462_113 : GEN_641;
  assign GEN_643 = 7'h72 == T_7300 ? T_10462_114 : GEN_642;
  assign GEN_644 = 7'h73 == T_7300 ? T_10462_115 : GEN_643;
  assign GEN_645 = 7'h74 == T_7300 ? T_10462_116 : GEN_644;
  assign GEN_646 = 7'h75 == T_7300 ? T_10462_117 : GEN_645;
  assign GEN_647 = 7'h76 == T_7300 ? T_10462_118 : GEN_646;
  assign GEN_648 = 7'h77 == T_7300 ? T_10462_119 : GEN_647;
  assign GEN_649 = 7'h78 == T_7300 ? T_10462_120 : GEN_648;
  assign GEN_650 = 7'h79 == T_7300 ? T_10462_121 : GEN_649;
  assign GEN_651 = 7'h7a == T_7300 ? T_10462_122 : GEN_650;
  assign GEN_652 = 7'h7b == T_7300 ? T_10462_123 : GEN_651;
  assign GEN_653 = 7'h7c == T_7300 ? T_10462_124 : GEN_652;
  assign GEN_654 = 7'h7d == T_7300 ? T_10462_125 : GEN_653;
  assign GEN_655 = 7'h7e == T_7300 ? T_10462_126 : GEN_654;
  assign GEN_656 = 7'h7f == T_7300 ? T_10462_127 : GEN_655;
  assign GEN_5 = GEN_783;
  assign GEN_657 = 7'h1 == T_7300 ? T_10725_1 : T_10725_0;
  assign GEN_658 = 7'h2 == T_7300 ? T_10725_2 : GEN_657;
  assign GEN_659 = 7'h3 == T_7300 ? T_10725_3 : GEN_658;
  assign GEN_660 = 7'h4 == T_7300 ? T_10725_4 : GEN_659;
  assign GEN_661 = 7'h5 == T_7300 ? T_10725_5 : GEN_660;
  assign GEN_662 = 7'h6 == T_7300 ? T_10725_6 : GEN_661;
  assign GEN_663 = 7'h7 == T_7300 ? T_10725_7 : GEN_662;
  assign GEN_664 = 7'h8 == T_7300 ? T_10725_8 : GEN_663;
  assign GEN_665 = 7'h9 == T_7300 ? T_10725_9 : GEN_664;
  assign GEN_666 = 7'ha == T_7300 ? T_10725_10 : GEN_665;
  assign GEN_667 = 7'hb == T_7300 ? T_10725_11 : GEN_666;
  assign GEN_668 = 7'hc == T_7300 ? T_10725_12 : GEN_667;
  assign GEN_669 = 7'hd == T_7300 ? T_10725_13 : GEN_668;
  assign GEN_670 = 7'he == T_7300 ? T_10725_14 : GEN_669;
  assign GEN_671 = 7'hf == T_7300 ? T_10725_15 : GEN_670;
  assign GEN_672 = 7'h10 == T_7300 ? T_10725_16 : GEN_671;
  assign GEN_673 = 7'h11 == T_7300 ? T_10725_17 : GEN_672;
  assign GEN_674 = 7'h12 == T_7300 ? T_10725_18 : GEN_673;
  assign GEN_675 = 7'h13 == T_7300 ? T_10725_19 : GEN_674;
  assign GEN_676 = 7'h14 == T_7300 ? T_10725_20 : GEN_675;
  assign GEN_677 = 7'h15 == T_7300 ? T_10725_21 : GEN_676;
  assign GEN_678 = 7'h16 == T_7300 ? T_10725_22 : GEN_677;
  assign GEN_679 = 7'h17 == T_7300 ? T_10725_23 : GEN_678;
  assign GEN_680 = 7'h18 == T_7300 ? T_10725_24 : GEN_679;
  assign GEN_681 = 7'h19 == T_7300 ? T_10725_25 : GEN_680;
  assign GEN_682 = 7'h1a == T_7300 ? T_10725_26 : GEN_681;
  assign GEN_683 = 7'h1b == T_7300 ? T_10725_27 : GEN_682;
  assign GEN_684 = 7'h1c == T_7300 ? T_10725_28 : GEN_683;
  assign GEN_685 = 7'h1d == T_7300 ? T_10725_29 : GEN_684;
  assign GEN_686 = 7'h1e == T_7300 ? T_10725_30 : GEN_685;
  assign GEN_687 = 7'h1f == T_7300 ? T_10725_31 : GEN_686;
  assign GEN_688 = 7'h20 == T_7300 ? T_10725_32 : GEN_687;
  assign GEN_689 = 7'h21 == T_7300 ? T_10725_33 : GEN_688;
  assign GEN_690 = 7'h22 == T_7300 ? T_10725_34 : GEN_689;
  assign GEN_691 = 7'h23 == T_7300 ? T_10725_35 : GEN_690;
  assign GEN_692 = 7'h24 == T_7300 ? T_10725_36 : GEN_691;
  assign GEN_693 = 7'h25 == T_7300 ? T_10725_37 : GEN_692;
  assign GEN_694 = 7'h26 == T_7300 ? T_10725_38 : GEN_693;
  assign GEN_695 = 7'h27 == T_7300 ? T_10725_39 : GEN_694;
  assign GEN_696 = 7'h28 == T_7300 ? T_10725_40 : GEN_695;
  assign GEN_697 = 7'h29 == T_7300 ? T_10725_41 : GEN_696;
  assign GEN_698 = 7'h2a == T_7300 ? T_10725_42 : GEN_697;
  assign GEN_699 = 7'h2b == T_7300 ? T_10725_43 : GEN_698;
  assign GEN_700 = 7'h2c == T_7300 ? T_10725_44 : GEN_699;
  assign GEN_701 = 7'h2d == T_7300 ? T_10725_45 : GEN_700;
  assign GEN_702 = 7'h2e == T_7300 ? T_10725_46 : GEN_701;
  assign GEN_703 = 7'h2f == T_7300 ? T_10725_47 : GEN_702;
  assign GEN_704 = 7'h30 == T_7300 ? T_10725_48 : GEN_703;
  assign GEN_705 = 7'h31 == T_7300 ? T_10725_49 : GEN_704;
  assign GEN_706 = 7'h32 == T_7300 ? T_10725_50 : GEN_705;
  assign GEN_707 = 7'h33 == T_7300 ? T_10725_51 : GEN_706;
  assign GEN_708 = 7'h34 == T_7300 ? T_10725_52 : GEN_707;
  assign GEN_709 = 7'h35 == T_7300 ? T_10725_53 : GEN_708;
  assign GEN_710 = 7'h36 == T_7300 ? T_10725_54 : GEN_709;
  assign GEN_711 = 7'h37 == T_7300 ? T_10725_55 : GEN_710;
  assign GEN_712 = 7'h38 == T_7300 ? T_10725_56 : GEN_711;
  assign GEN_713 = 7'h39 == T_7300 ? T_10725_57 : GEN_712;
  assign GEN_714 = 7'h3a == T_7300 ? T_10725_58 : GEN_713;
  assign GEN_715 = 7'h3b == T_7300 ? T_10725_59 : GEN_714;
  assign GEN_716 = 7'h3c == T_7300 ? T_10725_60 : GEN_715;
  assign GEN_717 = 7'h3d == T_7300 ? T_10725_61 : GEN_716;
  assign GEN_718 = 7'h3e == T_7300 ? T_10725_62 : GEN_717;
  assign GEN_719 = 7'h3f == T_7300 ? T_10725_63 : GEN_718;
  assign GEN_720 = 7'h40 == T_7300 ? T_10725_64 : GEN_719;
  assign GEN_721 = 7'h41 == T_7300 ? T_10725_65 : GEN_720;
  assign GEN_722 = 7'h42 == T_7300 ? T_10725_66 : GEN_721;
  assign GEN_723 = 7'h43 == T_7300 ? T_10725_67 : GEN_722;
  assign GEN_724 = 7'h44 == T_7300 ? T_10725_68 : GEN_723;
  assign GEN_725 = 7'h45 == T_7300 ? T_10725_69 : GEN_724;
  assign GEN_726 = 7'h46 == T_7300 ? T_10725_70 : GEN_725;
  assign GEN_727 = 7'h47 == T_7300 ? T_10725_71 : GEN_726;
  assign GEN_728 = 7'h48 == T_7300 ? T_10725_72 : GEN_727;
  assign GEN_729 = 7'h49 == T_7300 ? T_10725_73 : GEN_728;
  assign GEN_730 = 7'h4a == T_7300 ? T_10725_74 : GEN_729;
  assign GEN_731 = 7'h4b == T_7300 ? T_10725_75 : GEN_730;
  assign GEN_732 = 7'h4c == T_7300 ? T_10725_76 : GEN_731;
  assign GEN_733 = 7'h4d == T_7300 ? T_10725_77 : GEN_732;
  assign GEN_734 = 7'h4e == T_7300 ? T_10725_78 : GEN_733;
  assign GEN_735 = 7'h4f == T_7300 ? T_10725_79 : GEN_734;
  assign GEN_736 = 7'h50 == T_7300 ? T_10725_80 : GEN_735;
  assign GEN_737 = 7'h51 == T_7300 ? T_10725_81 : GEN_736;
  assign GEN_738 = 7'h52 == T_7300 ? T_10725_82 : GEN_737;
  assign GEN_739 = 7'h53 == T_7300 ? T_10725_83 : GEN_738;
  assign GEN_740 = 7'h54 == T_7300 ? T_10725_84 : GEN_739;
  assign GEN_741 = 7'h55 == T_7300 ? T_10725_85 : GEN_740;
  assign GEN_742 = 7'h56 == T_7300 ? T_10725_86 : GEN_741;
  assign GEN_743 = 7'h57 == T_7300 ? T_10725_87 : GEN_742;
  assign GEN_744 = 7'h58 == T_7300 ? T_10725_88 : GEN_743;
  assign GEN_745 = 7'h59 == T_7300 ? T_10725_89 : GEN_744;
  assign GEN_746 = 7'h5a == T_7300 ? T_10725_90 : GEN_745;
  assign GEN_747 = 7'h5b == T_7300 ? T_10725_91 : GEN_746;
  assign GEN_748 = 7'h5c == T_7300 ? T_10725_92 : GEN_747;
  assign GEN_749 = 7'h5d == T_7300 ? T_10725_93 : GEN_748;
  assign GEN_750 = 7'h5e == T_7300 ? T_10725_94 : GEN_749;
  assign GEN_751 = 7'h5f == T_7300 ? T_10725_95 : GEN_750;
  assign GEN_752 = 7'h60 == T_7300 ? T_10725_96 : GEN_751;
  assign GEN_753 = 7'h61 == T_7300 ? T_10725_97 : GEN_752;
  assign GEN_754 = 7'h62 == T_7300 ? T_10725_98 : GEN_753;
  assign GEN_755 = 7'h63 == T_7300 ? T_10725_99 : GEN_754;
  assign GEN_756 = 7'h64 == T_7300 ? T_10725_100 : GEN_755;
  assign GEN_757 = 7'h65 == T_7300 ? T_10725_101 : GEN_756;
  assign GEN_758 = 7'h66 == T_7300 ? T_10725_102 : GEN_757;
  assign GEN_759 = 7'h67 == T_7300 ? T_10725_103 : GEN_758;
  assign GEN_760 = 7'h68 == T_7300 ? T_10725_104 : GEN_759;
  assign GEN_761 = 7'h69 == T_7300 ? T_10725_105 : GEN_760;
  assign GEN_762 = 7'h6a == T_7300 ? T_10725_106 : GEN_761;
  assign GEN_763 = 7'h6b == T_7300 ? T_10725_107 : GEN_762;
  assign GEN_764 = 7'h6c == T_7300 ? T_10725_108 : GEN_763;
  assign GEN_765 = 7'h6d == T_7300 ? T_10725_109 : GEN_764;
  assign GEN_766 = 7'h6e == T_7300 ? T_10725_110 : GEN_765;
  assign GEN_767 = 7'h6f == T_7300 ? T_10725_111 : GEN_766;
  assign GEN_768 = 7'h70 == T_7300 ? T_10725_112 : GEN_767;
  assign GEN_769 = 7'h71 == T_7300 ? T_10725_113 : GEN_768;
  assign GEN_770 = 7'h72 == T_7300 ? T_10725_114 : GEN_769;
  assign GEN_771 = 7'h73 == T_7300 ? T_10725_115 : GEN_770;
  assign GEN_772 = 7'h74 == T_7300 ? T_10725_116 : GEN_771;
  assign GEN_773 = 7'h75 == T_7300 ? T_10725_117 : GEN_772;
  assign GEN_774 = 7'h76 == T_7300 ? T_10725_118 : GEN_773;
  assign GEN_775 = 7'h77 == T_7300 ? T_10725_119 : GEN_774;
  assign GEN_776 = 7'h78 == T_7300 ? T_10725_120 : GEN_775;
  assign GEN_777 = 7'h79 == T_7300 ? T_10725_121 : GEN_776;
  assign GEN_778 = 7'h7a == T_7300 ? T_10725_122 : GEN_777;
  assign GEN_779 = 7'h7b == T_7300 ? T_10725_123 : GEN_778;
  assign GEN_780 = 7'h7c == T_7300 ? T_10725_124 : GEN_779;
  assign GEN_781 = 7'h7d == T_7300 ? T_10725_125 : GEN_780;
  assign GEN_782 = 7'h7e == T_7300 ? T_10725_126 : GEN_781;
  assign GEN_783 = 7'h7f == T_7300 ? T_10725_127 : GEN_782;
  assign T_10858 = GEN_4 ? GEN_5 : 32'h0;
  assign T_10859 = T_992_bits_extra[9:8];
  assign T_10861 = T_992_bits_extra[7:3];
  assign T_10862 = T_992_bits_extra[2:0];
  assign T_10873_opcode = 3'h0;
  assign T_10873_param = 2'h0;
  assign T_10873_size = T_10862;
  assign T_10873_source = T_10861;
  assign T_10873_sink = 1'h0;
  assign T_10873_addr_lo = T_10859;
  assign T_10873_data = 32'h0;
  assign T_10873_error = 1'h0;

  always @(posedge clock) begin // Backup register no need to be reset
    if (T_3224) begin
      backupRegs_0 <= T_2505;
    end
    if (T_2984) begin
      backupRegs_1 <= T_2505;
    end
    if (T_3264) begin
      backupRegs_2 <= T_2505;
    end
    if (T_3784) begin
      backupRegs_3 <= T_2505;
    end
    if (T_4224) begin
      backupRegs_4 <= T_2505;
    end
    if (T_2664) begin
      backupRegs_5 <= T_2505;
    end
    if (T_2904) begin
      backupRegs_6 <= T_2505;
    end
    if (T_3624) begin
      backupRegs_7 <= T_2505;
    end
    if (T_4024) begin
      backupRegs_8 <= T_2505;
    end
    if (T_3104) begin
      backupRegs_9 <= T_2505;
    end
    if (T_2584) begin
      backupRegs_10 <= T_2505;
    end
    if (T_3984) begin
      backupRegs_11 <= T_2505;
    end
    if (T_3424) begin
      backupRegs_12 <= T_2505;
    end
    if (T_3304) begin
      backupRegs_13 <= T_2505;
    end
    if (T_2744) begin
      backupRegs_14 <= T_2505;
    end
    if (T_4384) begin
      backupRegs_15 <= T_2505;
    end
  end
endmodule
